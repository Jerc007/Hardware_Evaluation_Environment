
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity TP_instructions is
	port(
		instruction_pointer_in : in  integer;
		num_instructions_out   : out integer;
		instruction_out        : out std_logic_vector(31 downto 0)
	);
end TP_instructions;

architecture arch of TP_instructions is
	constant TP_INSTRUCTIONS : integer := 252;

begin
	num_instructions_out <= TP_INSTRUCTIONS;

	process(instruction_pointer_in)
	begin
		case instruction_pointer_in is
			when 0 => instruction_out <= x"d0800205";   -- 0000  LOP.AND.U16 R0H, R0H, c[0x1][0x0];    c[0x1][0x0] = 0x03ff
when 1 => instruction_out <= x"00400780";
when 2 => instruction_out <= x"a0000009";   -- 0008  I2I.U32.U16.C1 R2, R0L; 
when 3 => instruction_out <= x"040007d0";
when 4 => instruction_out <= x"a0000205";   -- 0010  I2I.U32.U16 R1, R0H; 
when 5 => instruction_out <= x"04000780";
when 6 => instruction_out <= x"a000f003";   -- 0018  SSY 0x78; 
when 7 => instruction_out <= x"00000000";
when 8 => instruction_out <= x"a0004e15";   -- 0020  I2I.U32.U16 R5, g [0x7].U16; 
when 9 => instruction_out <= x"04200780";
when 10 => instruction_out <= x"307c05fd";   -- 0028  ISET.S32.C0 o[0x7f], R2, R124, EQ; 
when 11 => instruction_out <= x"6c0087c8";
when 12 => instruction_out <= x"1000f003";   -- 0030  BRA C1.NEU, 0x78; 
when 13 => instruction_out <= x"00001680";
when 14 => instruction_out <= x"30040a01";   -- 0038  SHL R0, R5, 0x4; 
when 15 => instruction_out <= x"c4100780";
when 16 => instruction_out <= x"20000201";   -- 0040  IADD R0, R1, R0; 
when 17 => instruction_out <= x"04000780";
when 18 => instruction_out <= x"30020001";   -- 0048  SHL R0, R0, 0x2; 
when 19 => instruction_out <= x"c4100780";
when 20 => instruction_out <= x"2000c801";   -- 0050  IADD R0, g [0x4], R0; 
when 21 => instruction_out <= x"04200780";
when 22 => instruction_out <= x"20048001";   -- 0058  IADD32I R0, R0, 0x4; 
when 23 => instruction_out <= x"00000003";
when 24 => instruction_out <= x"d00e0001";   -- 0060  GLD.U32 R0, global14[R0]; 
when 25 => instruction_out <= x"80c00780";
when 26 => instruction_out <= x"00020205";   -- 0068  R2A A1, R1, 0x2; 
when 27 => instruction_out <= x"c0000780";
when 28 => instruction_out <= x"04001c01";   -- 0070  R2G.U32.U32 g[A1+0xe], R0; 
when 29 => instruction_out <= x"e4200780";
when 30 => instruction_out <= x"f0000001";   -- 0078  NOP.S; 
when 31 => instruction_out <= x"e0000002";
when 32 => instruction_out <= x"861ffe03";   -- 0080  BAR.ARV.WAIT b0, 0xfff; 
when 33 => instruction_out <= x"00000000";
when 34 => instruction_out <= x"3004d00d";   -- 0088  SHL R3, g [0x8], 0x4;  +-8
when 35 => instruction_out <= x"c4300780";
when 36 => instruction_out <= x"2101f001";   -- 0090  IADD32I R0, g [0x8], 0x1; +-8
when 37 => instruction_out <= x"00000003";
when 38 => instruction_out <= x"2010860d";   -- 0098  IADD32I R3, R3, 0x10; 
when 39 => instruction_out <= x"00000003";
when 40 => instruction_out <= x"40030010";   -- 00a0  IMUL32.U16.U16 R4, R0L, R1H;
when 41 => instruction_out <= x"400b0c18";   -- 00a4  IMUL32.U16.U16 R6, R3L, R5H;
when 42 => instruction_out <= x"60020211";   -- 00a8  IMAD.U16 R4, R0H, R1L, R4; 
when 43 => instruction_out <= x"00010780";
when 44 => instruction_out <= x"600a0e19";   -- 00b0  IMAD.U16 R6, R3H, R5L, R6; 
when 45 => instruction_out <= x"00018780";
when 46 => instruction_out <= x"30100811";   -- 00b8  SHL R4, R4, 0x10; 
when 47 => instruction_out <= x"c4100780";
when 48 => instruction_out <= x"30100c19";   -- 00c0  SHL R6, R6, 0x10; 
when 49 => instruction_out <= x"c4100780";
when 50 => instruction_out <= x"60020001";   -- 00c8  IMAD.U16 R0, R0L, R1L, R4; 
when 51 => instruction_out <= x"00010780";
when 52 => instruction_out <= x"600a0c0d";   -- 00d0  IMAD.U16 R3, R3L, R5L, R6; 
when 53 => instruction_out <= x"00018780";
when 54 => instruction_out <= x"20038000";   -- 00d8  IADD32 R0, R0, R3;
when 55 => instruction_out <= x"20008400";   -- 00dc  IADD32 R0, R2, R0;
when 56 => instruction_out <= x"2000d001";   -- 00e0  IADD R0, g [0x8], R0; +-8
when 57 => instruction_out <= x"04200780";
when 58 => instruction_out <= x"30020001";   -- 00e8  SHL R0, R0, 0x2; 
when 59 => instruction_out <= x"c4100780";
when 60 => instruction_out <= x"3004020d";   -- 00f0  SHL R3, R1, 0x4; 
when 61 => instruction_out <= x"c4100780";
when 62 => instruction_out <= x"2100ea18";   -- 00f8  IADD32 R6, g [0x5], R0;  +-5
when 63 => instruction_out <= x"2003840c";   -- 00fc  IADD32 R3, R2, R3;
when 64 => instruction_out <= x"20088c01";   -- 0100  IADD32I R0, R6, 0x8; 
when 65 => instruction_out <= x"00000003";
when 66 => instruction_out <= x"d00e0001";   -- 0108  GLD.U32 R0, global14[R0]; 
when 67 => instruction_out <= x"80c00780";
when 68 => instruction_out <= x"00020605";   -- 0110  R2A A1, R3, 0x2; 
when 69 => instruction_out <= x"c0000780";
when 70 => instruction_out <= x"04003c01";   -- 0118  R2G.U32.U32 g[A1+0x1e], R0; 
when 71 => instruction_out <= x"e4200780";
when 72 => instruction_out <= x"861ffe03";   -- 0120  BAR.ARV.WAIT b0, 0xfff; 
when 73 => instruction_out <= x"00000000";
when 74 => instruction_out <= x"00020209";   -- 0128  R2A A2, R1, 0x2; 
when 75 => instruction_out <= x"c0000780";
when 76 => instruction_out <= x"1400fc01";   -- 0130  MOV R0, g [A1+0x1e]; 
when 77 => instruction_out <= x"0423c780";
when 78 => instruction_out <= x"c800dc01";   -- 0138  FMUL R0, g [A2+0xe], R0; 
when 79 => instruction_out <= x"00200780";
when 80 => instruction_out <= x"04003c01";   -- 0140  R2G.U32.U32 g[A1+0x1e], R0; 
when 81 => instruction_out <= x"e4200780";
when 82 => instruction_out <= x"861ffe03";   -- 0148  BAR.ARV.WAIT b0, 0xfff; 
when 83 => instruction_out <= x"00000000";
when 84 => instruction_out <= x"10008001";   -- 0150  MVI R0, 0x3f800000; 
when 85 => instruction_out <= x"03f80003";
when 86 => instruction_out <= x"1001801d";   -- 0158  MVI R7, 0x1; 
when 87 => instruction_out <= x"00000003";
when 88 => instruction_out <= x"c0000001";   -- 0160  FMUL32I R0, R0, 0x3f800000; 
when 89 => instruction_out <= x"03f80003";
when 90 => instruction_out <= x"b0000001";   -- 0168  RRO R0, R0, EX2; 
when 91 => instruction_out <= x"c0004780";
when 92 => instruction_out <= x"90000001";   -- 0170  EX2 R0, R0; 
when 93 => instruction_out <= x"c0000780";
when 94 => instruction_out <= x"a000000d";   -- 0178  F2I.S32.F32.TRUNC R3, R0; 
when 95 => instruction_out <= x"8c064780";
when 96 => instruction_out <= x"10008200";   -- 0180  MOV32 R0, R1;
when 97 => instruction_out <= x"10008610";   -- 0184  MOV32 R4, R3;
when 98 => instruction_out <= x"20058003";   -- 0188  CAL.NOINC 0x2c0; 
when 99 => instruction_out <= x"00000000";
when 100 => instruction_out <= x"307c01fd";   -- 0190  ISET.S32.C1 o[0x7f], R0, R124, NE; 
when 101 => instruction_out <= x"6c0147d8";
when 102 => instruction_out <= x"a0040003";   -- 0198  SSY 0x200; 
when 103 => instruction_out <= x"00000000";
when 104 => instruction_out <= x"10040003";   -- 01a0  BRA C1.NE, 0x200; 
when 105 => instruction_out <= x"00001280";
when 106 => instruction_out <= x"301f0601";   -- 01a8  SHR.S32 R0, R3, 0x1f; 
when 107 => instruction_out <= x"ec100780";
when 108 => instruction_out <= x"d0810001";   -- 01b0  LOP.AND R0, R0, c[0x1][0x1];    c[0x1][0x1] = 0x10 or FFFFF
when 109 => instruction_out <= x"04400780";
when 110 => instruction_out <= x"20000001";   -- 01b8  IADD R0, R0, R3; 
when 111 => instruction_out <= x"0400c780";
when 112 => instruction_out <= x"30010001";   -- 01c0  SHR.S32 R0, R0, 0x1; 
when 113 => instruction_out <= x"ec100780";
when 114 => instruction_out <= x"20000201";   -- 01c8  IADD R0, R1, R0; 
when 115 => instruction_out <= x"04000780";
when 116 => instruction_out <= x"30040001";   -- 01d0  SHL R0, R0, 0x4; 
when 117 => instruction_out <= x"c4100780";
when 118 => instruction_out <= x"20000401";   -- 01d8  IADD R0, R2, R0; 
when 119 => instruction_out <= x"04000780";
when 120 => instruction_out <= x"00020009";   -- 01e0  R2A A2, R0, 0x2; 
when 121 => instruction_out <= x"c0000780";
when 122 => instruction_out <= x"1800fc01";   -- 01e8  MOV R0, g [A2+0x1e]; 
when 123 => instruction_out <= x"0423c780";
when 124 => instruction_out <= x"b400fc01";   -- 01f0  FADD R0, g [A1+0x1e], R0; 
when 125 => instruction_out <= x"00200780";
when 126 => instruction_out <= x"04003c01";   -- 01f8  R2G.U32.U32 g[A1+0x1e], R0; 
when 127 => instruction_out <= x"e4200780";
when 128 => instruction_out <= x"f0000001";   -- 0200  NOP.S; 
when 129 => instruction_out <= x"e0000002";
when 130 => instruction_out <= x"861ffe03";   -- 0208  BAR.ARV.WAIT b0, 0xfff; 
when 131 => instruction_out <= x"00000000";
when 132 => instruction_out <= x"20018e1d";   -- 0210  IADD32I R7, R7, 0x1; 
when 133 => instruction_out <= x"00000003";
when 134 => instruction_out <= x"a0000e01";   -- 0218  I2F.F32.S32 R0, R7; 
when 135 => instruction_out <= x"44014780";
when 136 => instruction_out <= x"b08201fd";   -- 0220  FSET.C1 o[0x7f], R0, c[0x1][0x2], LE; 	+-	c[0x1][0x2] = 4 but in float 0x40800000
when 137 => instruction_out <= x"6040c7d8";
when 138 => instruction_out <= x"1002c003";   -- 0228  BRA C1.NE, 0x160; 
when 139 => instruction_out <= x"00001280";
when 140 => instruction_out <= x"20088c0d";   -- 0230  IADD32I R3, R6, 0x8; 
when 141 => instruction_out <= x"00000003";
when 142 => instruction_out <= x"1400fc01";   -- 0238  MOV R0, g [A1+0x1e]; 
when 143 => instruction_out <= x"0423c780";
when 144 => instruction_out <= x"d00e0601";   -- 0240  GST.U32 global14[R3], R0; 
when 145 => instruction_out <= x"a0c00780";
when 146 => instruction_out <= x"861ffe03";   -- 0248  BAR.ARV.WAIT b0, 0xfff; 
when 147 => instruction_out <= x"00000000";
when 148 => instruction_out <= x"30000003";   -- 0250  RET C0.EQ; 
when 149 => instruction_out <= x"00000100";
when 150 => instruction_out <= x"1000d001";   -- 0258  MOV R0, g [0x8]; -8
when 151 => instruction_out <= x"0423c780";
when 152 => instruction_out <= x"4001140d";   -- 0260  IMUL.U16.U16 R3, R5L, R0H; 
when 153 => instruction_out <= x"00000780";
when 154 => instruction_out <= x"6000160d";   -- 0268  IMAD.U16 R3, R5H, R0L, R3; 
when 155 => instruction_out <= x"0000c780";
when 156 => instruction_out <= x"3010060d";   -- 0270  SHL R3, R3, 0x10; 
when 157 => instruction_out <= x"c4100780";
when 158 => instruction_out <= x"30040409";   -- 0278  SHL R2, R2, 0x4; 
when 159 => instruction_out <= x"c4100780";
when 160 => instruction_out <= x"60001401";   -- 0280  IMAD.U16 R0, R5L, R0L, R3; 
when 161 => instruction_out <= x"0000c780";
when 162 => instruction_out <= x"20028208";   -- 0288  IADD32 R2, R1, R2;
when 163 => instruction_out <= x"20018000";   -- 028c  IADD32 R0, R0, R1;
when 164 => instruction_out <= x"00020405";   -- 0290  R2A A1, R2, 0x2; 
when 165 => instruction_out <= x"c0000780";
when 166 => instruction_out <= x"30020005";   -- 0298  SHL R1, R0, 0x2; 
when 167 => instruction_out <= x"c4100780";
when 168 => instruction_out <= x"1400fc01";   -- 02a0  MOV R0, g [A1+0x1e]; 
when 169 => instruction_out <= x"0423c780";
when 170 => instruction_out <= x"2000cc05";   -- 02a8  IADD R1, g [0x6], R1; --6
when 171 => instruction_out <= x"04204780";
when 172 => instruction_out <= x"d00e0201";   -- 02b0  GST.U32 global14[R1], R0; 
when 173 => instruction_out <= x"a0c00780";
when 174 => instruction_out <= x"30000003";   -- 02b8  RET ; 
when 175 => instruction_out <= x"00000780";
when 176 => instruction_out <= x"a0000821";   -- 02c0  I2I.U32.S32 R8, |R4|; 
when 177 => instruction_out <= x"04114780";
when 178 => instruction_out <= x"a0001025";   -- 02c8  I2F.F32.U32 R9, R8; 
when 179 => instruction_out <= x"44004780";
when 180 => instruction_out <= x"a0000029";   -- 02d0  I2I.U32.S32 R10, |R0|; 
when 181 => instruction_out <= x"04114780";
when 182 => instruction_out <= x"9000122d";   -- 02d8  RCP R11, R9; 
when 183 => instruction_out <= x"00000780";
when 184 => instruction_out <= x"a0001425";   -- 02e0  I2F.F32.U32.TRUNC R9, R10; 
when 185 => instruction_out <= x"44064780";
when 186 => instruction_out <= x"203e962d";   -- 02e8  IADD32I R11, R11, 0xfffffffe; 
when 187 => instruction_out <= x"0fffffff";
when 188 => instruction_out <= x"c00b1225";   -- 02f0  FMUL.TRUNC.C1 R9, R9, R11; 
when 189 => instruction_out <= x"0000c7d0";
when 190 => instruction_out <= x"a0001225";   -- 02f8  F2I.U32.F32.TRUNC R9, R9; 
when 191 => instruction_out <= x"84064780";
when 192 => instruction_out <= x"40132031";   -- 0300  IMUL.U16.U16 R12, R8L, R9H; 
when 193 => instruction_out <= x"00000780";
when 194 => instruction_out <= x"60122231";   -- 0308  IMAD.U16 R12, R8H, R9L, R12; 
when 195 => instruction_out <= x"00030780";
when 196 => instruction_out <= x"30101831";   -- 0310  SHL R12, R12, 0x10; 
when 197 => instruction_out <= x"c4100780";
when 198 => instruction_out <= x"60122031";   -- 0318  IMAD.U16 R12, R8L, R9L, R12; 
when 199 => instruction_out <= x"00030780";
when 200 => instruction_out <= x"20401431";   -- 0320  IADD R12, R10, -R12; 
when 201 => instruction_out <= x"04030780";
when 202 => instruction_out <= x"a0001831";   -- 0328  I2F.F32.U32.TRUNC R12, R12; 
when 203 => instruction_out <= x"44064780";
when 204 => instruction_out <= x"c00b182d";   -- 0330  FMUL.TRUNC.C1 R11, R12, R11; 
when 205 => instruction_out <= x"0000c7d0";
when 206 => instruction_out <= x"a000162d";   -- 0338  F2I.U32.F32.TRUNC R11, R11; 
when 207 => instruction_out <= x"84064780";
when 208 => instruction_out <= x"20001225";   -- 0340  IADD R9, R9, R11; 
when 209 => instruction_out <= x"0402c780";
when 210 => instruction_out <= x"4010262d";   -- 0348  IMUL.U16.U16 R11, R9H, R8L; 
when 211 => instruction_out <= x"00000780";
when 212 => instruction_out <= x"6011242d";   -- 0350  IMAD.U16 R11, R9L, R8H, R11; 
when 213 => instruction_out <= x"0002c780";
when 214 => instruction_out <= x"3010162d";   -- 0358  SHL R11, R11, 0x10; 
when 215 => instruction_out <= x"c4100780";
when 216 => instruction_out <= x"6010242d";   -- 0360  IMAD.U16 R11, R9L, R8L, R11; 
when 217 => instruction_out <= x"0002c780";
when 218 => instruction_out <= x"3000162d";   -- 0368  IADD R11, -R11, R10; 
when 219 => instruction_out <= x"04028780";
when 220 => instruction_out <= x"300b102d";   -- 0370  ISET R11, R8, R11, LE; 
when 221 => instruction_out <= x"6400c780";
when 222 => instruction_out <= x"30001625";   -- 0378  IADD R9, -R11, R9; 
when 223 => instruction_out <= x"04024780";
when 224 => instruction_out <= x"4010262d";   -- 0380  IMUL.U16.U16 R11, R9H, R8L; 
when 225 => instruction_out <= x"00000780";
when 226 => instruction_out <= x"6011242d";   -- 0388  IMAD.U16 R11, R9L, R8H, R11; 
when 227 => instruction_out <= x"0002c780";
when 228 => instruction_out <= x"3010162d";   -- 0390  SHL R11, R11, 0x10; 
when 229 => instruction_out <= x"c4100780";
when 230 => instruction_out <= x"60102421";   -- 0398  IMAD.U16 R8, R9L, R8L, R11; 
when 231 => instruction_out <= x"0002c780";
when 232 => instruction_out <= x"301f0001";   -- 03a0  SHR R0, R0, 0x1f; 
when 233 => instruction_out <= x"e4100780";
when 234 => instruction_out <= x"30001025";   -- 03a8  IADD R9, -R8, R10; 
when 235 => instruction_out <= x"04028780";
when 236 => instruction_out <= x"a0000021";   -- 03b0  I2I.S32.S32 R8, -R0; 
when 237 => instruction_out <= x"2c014780";
when 238 => instruction_out <= x"d0091021";   -- 03b8  LOP.XOR R8, R8, R9; 
when 239 => instruction_out <= x"04008780";
when 240 => instruction_out <= x"307c09fd";   -- 03c0  ISET.S32.C1 o[0x7f], R4, R124, NE; 
when 241 => instruction_out <= x"6c0147d8";
when 242 => instruction_out <= x"20000001";   -- 03c8  IADD R0, R0, R8; 
when 243 => instruction_out <= x"04020780";
when 244 => instruction_out <= x"d0040001";   -- 03d0  LOP.PASS_B R0 (C1.EQU), R0, ~R4; 
when 245 => instruction_out <= x"0402d500";
when 246 => instruction_out <= x"30000003";   -- 03d8  RET C1; 
when 247 => instruction_out <= x"00001780";
when 248 => instruction_out <= x"f0000001";   -- 03e0  NOP; 
when 249 => instruction_out <= x"e0000001";
when 250 => instruction_out <= x"30000003";   -- RET ;
when 251 => instruction_out <= x"00000780";

			when others => null;
		end case;
	end process;

end arch;
