
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity TP_instructions is
	port(
		instruction_pointer_in : in  integer;
		num_instructions_out   : out integer;
		instruction_out        : out std_logic_vector(31 downto 0)
	);
end TP_instructions;

architecture arch of TP_instructions is
	constant TP_INSTRUCTIONS : integer := 336;

begin
	num_instructions_out <= TP_INSTRUCTIONS;

	process(instruction_pointer_in)
	begin
		case instruction_pointer_in is
			when 0 => instruction_out <= x"a0004e09";   -- 0000  I2I.U32.U16 R2, g [0x7].U16; 
when 1 => instruction_out <= x"04200780";
when 2 => instruction_out <= x"1000ce05";   -- 0008  MOV R1, g [0x7]; 
when 3 => instruction_out <= x"0423c780";
when 4 => instruction_out <= x"4003080d";   -- 0010  IMUL.U16.U16 R3, R2L, R1H; 
when 5 => instruction_out <= x"00000780";
when 6 => instruction_out <= x"60020a0d";   -- 0018  IMAD.U16 R3, R2H, R1L, R3; 
when 7 => instruction_out <= x"0000c780";
when 8 => instruction_out <= x"3010060d";   -- 0020  SHL R3, R3, 0x10; 
when 9 => instruction_out <= x"c4100780";
when 10 => instruction_out <= x"60020805";   -- 0028  IMAD.U16 R1, R2L, R1L, R3; 
when 11 => instruction_out <= x"0000c780";
when 12 => instruction_out <= x"30050219";   -- 0030  SHL R6, R1, 0x5; 
when 13 => instruction_out <= x"c4100780";
when 14 => instruction_out <= x"2000ce05";   -- 0038  IADD R1, g [0x7], R6; 
when 15 => instruction_out <= x"04218780";
when 16 => instruction_out <= x"203f821d";   -- 0040  IADD32I R7, R1, 0xffffffff; 
when 17 => instruction_out <= x"0fffffff";
when 18 => instruction_out <= x"a0004c0d";   -- 0048  I2I.U32.U16 R3, g [0x6].U16; 
when 19 => instruction_out <= x"04200780";
when 20 => instruction_out <= x"d0800205";   -- 0050  LOP.AND.U16 R0H, R0H, c[0x1][0x0]; 
when 21 => instruction_out <= x"00400780";
when 22 => instruction_out <= x"30060ffd";   -- 0058  ISET.S32.C0 o[0x7f], R7, R6, LT; 
when 23 => instruction_out <= x"6c0047c8";
when 24 => instruction_out <= x"30050621";   -- 0060  SHL R8, R3, 0x5; 
when 25 => instruction_out <= x"c4100780";
when 26 => instruction_out <= x"a0000011";   -- 0068  I2I.U32.U16 R4, R0L; 
when 27 => instruction_out <= x"04000780";
when 28 => instruction_out <= x"a0000215";   -- 0070  I2I.U32.U16 R5, R0H; 
when 29 => instruction_out <= x"04000780";
when 30 => instruction_out <= x"10096003";   -- 0078  BRA C0.NE, 0x4b0; 
when 31 => instruction_out <= x"00000280";
when 32 => instruction_out <= x"1100f004";   -- 0080  MOV32 R1, g [0x8];
when 33 => instruction_out <= x"1100ee00";   -- 0084  MOV32 R0, g [0x7];
when 34 => instruction_out <= x"4003142c";   -- 0088  IMUL32.U16.U16 R11, R5L, R1H;
when 35 => instruction_out <= x"40011424";   -- 008c  IMUL32.U16.U16 R9, R5L, R0H;
when 36 => instruction_out <= x"30050a29";   -- 0090  SHL R10, R5, 0x5; 
when 37 => instruction_out <= x"c4100780";
when 38 => instruction_out <= x"60021631";   -- 0098  IMAD.U16 R12, R5H, R1L, R11; 
when 39 => instruction_out <= x"0002c780";
when 40 => instruction_out <= x"60001625";   -- 00a0  IMAD.U16 R9, R5H, R0L, R9; 
when 41 => instruction_out <= x"00024780";
when 42 => instruction_out <= x"30070a2d";   -- 00a8  SHL R11, R5, 0x7; 
when 43 => instruction_out <= x"c4100780";
when 44 => instruction_out <= x"20000829";   -- 00b0  IADD R10, R4, R10; 
when 45 => instruction_out <= x"04028780";
when 46 => instruction_out <= x"30101831";   -- 00b8  SHL R12, R12, 0x10; 
when 47 => instruction_out <= x"c4100780";
when 48 => instruction_out <= x"30101225";   -- 00c0  SHL R9, R9, 0x10; 
when 49 => instruction_out <= x"c4100780";
when 50 => instruction_out <= x"2030962d";   -- 00c8  IADD32I R11, R11, 0x30; 
when 51 => instruction_out <= x"00000003";
when 52 => instruction_out <= x"00021405";   -- 00d0  R2A A1, R10, 0x2; 
when 53 => instruction_out <= x"c0000780";
when 54 => instruction_out <= x"60021405";   -- 00d8  IMAD.U16 R1, R5L, R1L, R12; 
when 55 => instruction_out <= x"00030780";
when 56 => instruction_out <= x"60001401";   -- 00e0  IMAD.U16 R0, R5L, R0L, R9; 
when 57 => instruction_out <= x"00024780";
when 58 => instruction_out <= x"00001609";   -- 00e8  R2A A2, R11; 
when 59 => instruction_out <= x"c0000780";
when 60 => instruction_out <= x"200c8825";   -- 00f0  IADD32I R9, R4, 0x40c; 
when 61 => instruction_out <= x"00000043";
when 62 => instruction_out <= x"20088220";   -- 00f8  IADD32 R8, R1, R8;
when 63 => instruction_out <= x"20068014";   -- 00fc  IADD32 R5, R0, R6;
when 64 => instruction_out <= x"20000001";   -- 0100  IADD R0, R0, R7; 
when 65 => instruction_out <= x"0401c780";
when 66 => instruction_out <= x"0002120d";   -- 0108  R2A A3, R9, 0x2; 
when 67 => instruction_out <= x"c0000780";
when 68 => instruction_out <= x"20088818";   -- 0110  IADD32 R6, R4, R8;
when 69 => instruction_out <= x"20058820";   -- 0114  IADD32 R8, R4, R5;
when 70 => instruction_out <= x"a0094003";   -- 0118  SSY 0x4a0; 
when 71 => instruction_out <= x"00000000";
when 72 => instruction_out <= x"3007d01d";   -- 0120  SHL R7, g [0x8], 0x7; 
when 73 => instruction_out <= x"c4300780";
when 74 => instruction_out <= x"30020c19";   -- 0128  SHL R6, R6, 0x2; 
when 75 => instruction_out <= x"c4100780";
when 76 => instruction_out <= x"30021015";   -- 0130  SHL R5, R8, 0x2; 
when 77 => instruction_out <= x"c4100780";
when 78 => instruction_out <= x"1000f829";   -- 0138  MOV R10, R124; 
when 79 => instruction_out <= x"0403c780";
when 80 => instruction_out <= x"20008824";   -- 0140  IADD32 R9, R4, R0;
when 81 => instruction_out <= x"2106ec18";   -- 0144  IADD32 R6, g [0x6], R6;
when 82 => instruction_out <= x"2000ca15";   -- 0148  IADD R5, g [0x5], R5; 
when 83 => instruction_out <= x"04214780";
when 84 => instruction_out <= x"d00e0a2d";   -- 0150  GLD.U32 R11, global14[R5]; 
when 85 => instruction_out <= x"80c00780";
when 86 => instruction_out <= x"d00e0c01";   -- 0158  GLD.U32 R0, global14[R6]; 
when 87 => instruction_out <= x"80c00780";
when 88 => instruction_out <= x"04001801";   -- 0160  R2G.U32.U32 g[A1+0xc], R11; 
when 89 => instruction_out <= x"e422c780";
when 90 => instruction_out <= x"04081801";   -- 0168  R2G.U32.U32 g[A1+0x40c], R0; 
when 91 => instruction_out <= x"e4200780";
when 92 => instruction_out <= x"861ffe03";   -- 0170  BAR.ARV.WAIT b0, 0xfff; 
when 93 => instruction_out <= x"00000000";
when 94 => instruction_out <= x"1c00c001";   -- 0178  MOV R0, g [A3+0x0]; 
when 95 => instruction_out <= x"0423c780";
when 96 => instruction_out <= x"dc010011";   -- 0180  ADA A4, A3, 0x80; 
when 97 => instruction_out <= x"20000780";
when 98 => instruction_out <= x"e800c029";   -- 0188  FMAD R10, g [A2+0x0], R0, R10; 
when 99 => instruction_out <= x"00228780";
when 100 => instruction_out <= x"1000c001";   -- 0190  MOV R0, g [A4+0x0]; 
when 101 => instruction_out <= x"0423c784";
when 102 => instruction_out <= x"dc020011";   -- 0198  ADA A4, A3, 0x100; 
when 103 => instruction_out <= x"20000780";
when 104 => instruction_out <= x"e800c229";   -- 01a0  FMAD R10, g [A2+0x1], R0, R10; 
when 105 => instruction_out <= x"00228780";
when 106 => instruction_out <= x"1000c001";   -- 01a8  MOV R0, g [A4+0x0]; 
when 107 => instruction_out <= x"0423c784";
when 108 => instruction_out <= x"dc030011";   -- 01b0  ADA A4, A3, 0x180; 
when 109 => instruction_out <= x"20000780";
when 110 => instruction_out <= x"e800c429";   -- 01b8  FMAD R10, g [A2+0x2], R0, R10; 
when 111 => instruction_out <= x"00228780";
when 112 => instruction_out <= x"1000c001";   -- 01c0  MOV R0, g [A4+0x0]; 
when 113 => instruction_out <= x"0423c784";
when 114 => instruction_out <= x"dc040011";   -- 01c8  ADA A4, A3, 0x200; 
when 115 => instruction_out <= x"20000780";
when 116 => instruction_out <= x"e800c629";   -- 01d0  FMAD R10, g [A2+0x3], R0, R10; 
when 117 => instruction_out <= x"00228780";
when 118 => instruction_out <= x"1000c001";   -- 01d8  MOV R0, g [A4+0x0]; 
when 119 => instruction_out <= x"0423c784";
when 120 => instruction_out <= x"dc050011";   -- 01e0  ADA A4, A3, 0x280; 
when 121 => instruction_out <= x"20000780";
when 122 => instruction_out <= x"e800c829";   -- 01e8  FMAD R10, g [A2+0x4], R0, R10; 
when 123 => instruction_out <= x"00228780";
when 124 => instruction_out <= x"1000c001";   -- 01f0  MOV R0, g [A4+0x0]; 
when 125 => instruction_out <= x"0423c784";
when 126 => instruction_out <= x"dc060011";   -- 01f8  ADA A4, A3, 0x300; 
when 127 => instruction_out <= x"20000780";
when 128 => instruction_out <= x"e800ca29";   -- 0200  FMAD R10, g [A2+0x5], R0, R10; 
when 129 => instruction_out <= x"00228780";
when 130 => instruction_out <= x"1000c001";   -- 0208  MOV R0, g [A4+0x0]; 
when 131 => instruction_out <= x"0423c784";
when 132 => instruction_out <= x"dc070011";   -- 0210  ADA A4, A3, 0x380; 
when 133 => instruction_out <= x"20000780";
when 134 => instruction_out <= x"e800cc29";   -- 0218  FMAD R10, g [A2+0x6], R0, R10; 
when 135 => instruction_out <= x"00228780";
when 136 => instruction_out <= x"1000c001";   -- 0220  MOV R0, g [A4+0x0]; 
when 137 => instruction_out <= x"0423c784";
when 138 => instruction_out <= x"dc080011";   -- 0228  ADA A4, A3, 0x400; 
when 139 => instruction_out <= x"20000780";
when 140 => instruction_out <= x"e800ce29";   -- 0230  FMAD R10, g [A2+0x7], R0, R10; 
when 141 => instruction_out <= x"00228780";
when 142 => instruction_out <= x"1000c001";   -- 0238  MOV R0, g [A4+0x0]; 
when 143 => instruction_out <= x"0423c784";
when 144 => instruction_out <= x"dc090011";   -- 0240  ADA A4, A3, 0x480; 
when 145 => instruction_out <= x"20000780";
when 146 => instruction_out <= x"e800d029";   -- 0248  FMAD R10, g [A2+0x8], R0, R10; 
when 147 => instruction_out <= x"00228780";
when 148 => instruction_out <= x"1000c001";   -- 0250  MOV R0, g [A4+0x0]; 
when 149 => instruction_out <= x"0423c784";
when 150 => instruction_out <= x"dc0a0011";   -- 0258  ADA A4, A3, 0x500; 
when 151 => instruction_out <= x"20000780";
when 152 => instruction_out <= x"e800d229";   -- 0260  FMAD R10, g [A2+0x9], R0, R10; 
when 153 => instruction_out <= x"00228780";
when 154 => instruction_out <= x"1000c001";   -- 0268  MOV R0, g [A4+0x0]; 
when 155 => instruction_out <= x"0423c784";
when 156 => instruction_out <= x"dc0b0011";   -- 0270  ADA A4, A3, 0x580; 
when 157 => instruction_out <= x"20000780";
when 158 => instruction_out <= x"e800d429";   -- 0278  FMAD R10, g [A2+0xa], R0, R10; 
when 159 => instruction_out <= x"00228780";
when 160 => instruction_out <= x"1000c001";   -- 0280  MOV R0, g [A4+0x0]; 
when 161 => instruction_out <= x"0423c784";
when 162 => instruction_out <= x"dc0c0011";   -- 0288  ADA A4, A3, 0x600; 
when 163 => instruction_out <= x"20000780";
when 164 => instruction_out <= x"e800d629";   -- 0290  FMAD R10, g [A2+0xb], R0, R10; 
when 165 => instruction_out <= x"00228780";
when 166 => instruction_out <= x"1000c001";   -- 0298  MOV R0, g [A4+0x0]; 
when 167 => instruction_out <= x"0423c784";
when 168 => instruction_out <= x"dc0d0011";   -- 02a0  ADA A4, A3, 0x680; 
when 169 => instruction_out <= x"20000780";
when 170 => instruction_out <= x"e800d829";   -- 02a8  FMAD R10, g [A2+0xc], R0, R10; 
when 171 => instruction_out <= x"00228780";
when 172 => instruction_out <= x"1000c001";   -- 02b0  MOV R0, g [A4+0x0]; 
when 173 => instruction_out <= x"0423c784";
when 174 => instruction_out <= x"dc0e0011";   -- 02b8  ADA A4, A3, 0x700; 
when 175 => instruction_out <= x"20000780";
when 176 => instruction_out <= x"e800da29";   -- 02c0  FMAD R10, g [A2+0xd], R0, R10; 
when 177 => instruction_out <= x"00228780";
when 178 => instruction_out <= x"1000c001";   -- 02c8  MOV R0, g [A4+0x0]; 
when 179 => instruction_out <= x"0423c784";
when 180 => instruction_out <= x"dc0f0011";   -- 02d0  ADA A4, A3, 0x780; 
when 181 => instruction_out <= x"20000780";
when 182 => instruction_out <= x"e800dc29";   -- 02d8  FMAD R10, g [A2+0xe], R0, R10; 
when 183 => instruction_out <= x"00228780";
when 184 => instruction_out <= x"1000c001";   -- 02e0  MOV R0, g [A4+0x0]; 
when 185 => instruction_out <= x"0423c784";
when 186 => instruction_out <= x"dc100011";   -- 02e8  ADA A4, A3, 0x800; 
when 187 => instruction_out <= x"20000780";
when 188 => instruction_out <= x"e800de29";   -- 02f0  FMAD R10, g [A2+0xf], R0, R10; 
when 189 => instruction_out <= x"00228780";
when 190 => instruction_out <= x"1000c001";   -- 02f8  MOV R0, g [A4+0x0]; 
when 191 => instruction_out <= x"0423c784";
when 192 => instruction_out <= x"dc110011";   -- 0300  ADA A4, A3, 0x880; 
when 193 => instruction_out <= x"20000780";
when 194 => instruction_out <= x"e800e029";   -- 0308  FMAD R10, g [A2+0x10], R0, R10; 
when 195 => instruction_out <= x"00228780";
when 196 => instruction_out <= x"1000c001";   -- 0310  MOV R0, g [A4+0x0]; 
when 197 => instruction_out <= x"0423c784";
when 198 => instruction_out <= x"dc120011";   -- 0318  ADA A4, A3, 0x900; 
when 199 => instruction_out <= x"20000780";
when 200 => instruction_out <= x"e800e229";   -- 0320  FMAD R10, g [A2+0x11], R0, R10; 
when 201 => instruction_out <= x"00228780";
when 202 => instruction_out <= x"1000c001";   -- 0328  MOV R0, g [A4+0x0]; 
when 203 => instruction_out <= x"0423c784";
when 204 => instruction_out <= x"dc130011";   -- 0330  ADA A4, A3, 0x980; 
when 205 => instruction_out <= x"20000780";
when 206 => instruction_out <= x"e800e429";   -- 0338  FMAD R10, g [A2+0x12], R0, R10; 
when 207 => instruction_out <= x"00228780";
when 208 => instruction_out <= x"1000c001";   -- 0340  MOV R0, g [A4+0x0]; 
when 209 => instruction_out <= x"0423c784";
when 210 => instruction_out <= x"dc140011";   -- 0348  ADA A4, A3, 0xa00; 
when 211 => instruction_out <= x"20000780";
when 212 => instruction_out <= x"e800e629";   -- 0350  FMAD R10, g [A2+0x13], R0, R10; 
when 213 => instruction_out <= x"00228780";
when 214 => instruction_out <= x"1000c001";   -- 0358  MOV R0, g [A4+0x0]; 
when 215 => instruction_out <= x"0423c784";
when 216 => instruction_out <= x"dc150011";   -- 0360  ADA A4, A3, 0xa80; 
when 217 => instruction_out <= x"20000780";
when 218 => instruction_out <= x"e800e829";   -- 0368  FMAD R10, g [A2+0x14], R0, R10; 
when 219 => instruction_out <= x"00228780";
when 220 => instruction_out <= x"1000c001";   -- 0370  MOV R0, g [A4+0x0]; 
when 221 => instruction_out <= x"0423c784";
when 222 => instruction_out <= x"dc160011";   -- 0378  ADA A4, A3, 0xb00; 
when 223 => instruction_out <= x"20000780";
when 224 => instruction_out <= x"e800ea29";   -- 0380  FMAD R10, g [A2+0x15], R0, R10; 
when 225 => instruction_out <= x"00228780";
when 226 => instruction_out <= x"1000c001";   -- 0388  MOV R0, g [A4+0x0]; 
when 227 => instruction_out <= x"0423c784";
when 228 => instruction_out <= x"dc170011";   -- 0390  ADA A4, A3, 0xb80; 
when 229 => instruction_out <= x"20000780";
when 230 => instruction_out <= x"e800ec29";   -- 0398  FMAD R10, g [A2+0x16], R0, R10; 
when 231 => instruction_out <= x"00228780";
when 232 => instruction_out <= x"1000c001";   -- 03a0  MOV R0, g [A4+0x0]; 
when 233 => instruction_out <= x"0423c784";
when 234 => instruction_out <= x"dc180011";   -- 03a8  ADA A4, A3, 0xc00; 
when 235 => instruction_out <= x"20000780";
when 236 => instruction_out <= x"e800ee29";   -- 03b0  FMAD R10, g [A2+0x17], R0, R10; 
when 237 => instruction_out <= x"00228780";
when 238 => instruction_out <= x"1000c001";   -- 03b8  MOV R0, g [A4+0x0]; 
when 239 => instruction_out <= x"0423c784";
when 240 => instruction_out <= x"dc190011";   -- 03c0  ADA A4, A3, 0xc80; 
when 241 => instruction_out <= x"20000780";
when 242 => instruction_out <= x"e800f029";   -- 03c8  FMAD R10, g [A2+0x18], R0, R10; 
when 243 => instruction_out <= x"00228780";
when 244 => instruction_out <= x"1000c001";   -- 03d0  MOV R0, g [A4+0x0]; 
when 245 => instruction_out <= x"0423c784";
when 246 => instruction_out <= x"dc1a0011";   -- 03d8  ADA A4, A3, 0xd00; 
when 247 => instruction_out <= x"20000780";
when 248 => instruction_out <= x"e800f229";   -- 03e0  FMAD R10, g [A2+0x19], R0, R10; 
when 249 => instruction_out <= x"00228780";
when 250 => instruction_out <= x"1000c001";   -- 03e8  MOV R0, g [A4+0x0]; 
when 251 => instruction_out <= x"0423c784";
when 252 => instruction_out <= x"dc1b0011";   -- 03f0  ADA A4, A3, 0xd80; 
when 253 => instruction_out <= x"20000780";
when 254 => instruction_out <= x"e800f429";   -- 03f8  FMAD R10, g [A2+0x1a], R0, R10; 
when 255 => instruction_out <= x"00228780";
when 256 => instruction_out <= x"1000c001";   -- 0400  MOV R0, g [A4+0x0]; 
when 257 => instruction_out <= x"0423c784";
when 258 => instruction_out <= x"dc1c0011";   -- 0408  ADA A4, A3, 0xe00; 
when 259 => instruction_out <= x"20000780";
when 260 => instruction_out <= x"e800f629";   -- 0410  FMAD R10, g [A2+0x1b], R0, R10; 
when 261 => instruction_out <= x"00228780";
when 262 => instruction_out <= x"1000c001";   -- 0418  MOV R0, g [A4+0x0]; 
when 263 => instruction_out <= x"0423c784";
when 264 => instruction_out <= x"dc1d0011";   -- 0420  ADA A4, A3, 0xe80; 
when 265 => instruction_out <= x"20000780";
when 266 => instruction_out <= x"e800f829";   -- 0428  FMAD R10, g [A2+0x1c], R0, R10; 
when 267 => instruction_out <= x"00228780";
when 268 => instruction_out <= x"1000c001";   -- 0430  MOV R0, g [A4+0x0]; 
when 269 => instruction_out <= x"0423c784";
when 270 => instruction_out <= x"dc1e0011";   -- 0438  ADA A4, A3, 0xf00; 
when 271 => instruction_out <= x"20000780";
when 272 => instruction_out <= x"e800fa29";   -- 0440  FMAD R10, g [A2+0x1d], R0, R10; 
when 273 => instruction_out <= x"00228780";
when 274 => instruction_out <= x"1000c001";   -- 0448  MOV R0, g [A4+0x0]; 
when 275 => instruction_out <= x"0423c784";
when 276 => instruction_out <= x"dc1f0011";   -- 0450  ADA A4, A3, 0xf80; 
when 277 => instruction_out <= x"20000780";
when 278 => instruction_out <= x"e800fc29";   -- 0458  FMAD R10, g [A2+0x1e], R0, R10; 
when 279 => instruction_out <= x"00228780";
when 280 => instruction_out <= x"1000c001";   -- 0460  MOV R0, g [A4+0x0]; 
when 281 => instruction_out <= x"0423c784";
when 282 => instruction_out <= x"e800fe29";   -- 0468  FMAD R10, g [A2+0x1f], R0, R10; 
when 283 => instruction_out <= x"00228780";
when 284 => instruction_out <= x"861ffe03";   -- 0470  BAR.ARV.WAIT b0, 0xfff; 
when 285 => instruction_out <= x"00000000";
when 286 => instruction_out <= x"20209021";   -- 0478  IADD32I R8, R8, 0x20; 
when 287 => instruction_out <= x"00000003";
when 288 => instruction_out <= x"300911fd";   -- 0480  ISET.S32.C0 o[0x7f], R8, R9, LE; 
when 289 => instruction_out <= x"6c00c7c8";
when 290 => instruction_out <= x"20008a15";   -- 0488  IADD32I R5, R5, 0x80; 
when 291 => instruction_out <= x"0000000b";
when 292 => instruction_out <= x"20000e19";   -- 0490  IADD R6, R7, R6; 
when 293 => instruction_out <= x"04018780";
when 294 => instruction_out <= x"1002a003";   -- 0498  BRA C0.NE, 0x150; 
when 295 => instruction_out <= x"00000280";
when 296 => instruction_out <= x"f0000001";   -- 04a0  NOP.S; 
when 297 => instruction_out <= x"e0000002";
when 298 => instruction_out <= x"1009c003";   -- 04a8  BRA  0x4e0; 
when 299 => instruction_out <= x"00000780";
when 300 => instruction_out <= x"1000d001";   -- 04b0  MOV R0, g [0x8]; 
when 301 => instruction_out <= x"0423c780";
when 302 => instruction_out <= x"40011405";   -- 04b8  IMUL.U16.U16 R1, R5L, R0H; 
when 303 => instruction_out <= x"00000780";
when 304 => instruction_out <= x"60001605";   -- 04c0  IMAD.U16 R1, R5H, R0L, R1; 
when 305 => instruction_out <= x"00004780";
when 306 => instruction_out <= x"30100205";   -- 04c8  SHL R1, R1, 0x10; 
when 307 => instruction_out <= x"c4100780";
when 308 => instruction_out <= x"60001405";   -- 04d0  IMAD.U16 R1, R5L, R0L, R1; 
when 309 => instruction_out <= x"00004780";
when 310 => instruction_out <= x"1000f829";   -- 04d8  MOV R10, R124; 
when 311 => instruction_out <= x"0403c780";
when 312 => instruction_out <= x"1000d001";   -- 04e0  MOV R0, g [0x8]; 
when 313 => instruction_out <= x"0423c780";
when 314 => instruction_out <= x"40050015";   -- 04e8  IMUL.U16.U16 R5, R0L, R2H; 
when 315 => instruction_out <= x"00000780";
when 316 => instruction_out <= x"60040215";   -- 04f0  IMAD.U16 R5, R0H, R2L, R5; 
when 317 => instruction_out <= x"00014780";
when 318 => instruction_out <= x"30100a15";   -- 04f8  SHL R5, R5, 0x10; 
when 319 => instruction_out <= x"c4100780";
when 320 => instruction_out <= x"60040001";   -- 0500  IMAD.U16 R0, R0L, R2L, R5; 
when 321 => instruction_out <= x"00014780";
when 322 => instruction_out <= x"20000001";   -- 0508  IADD R0, R0, R3; 
when 323 => instruction_out <= x"0400c780";
when 324 => instruction_out <= x"30050001";   -- 0510  SHL R0, R0, 0x5; 
when 325 => instruction_out <= x"c4100780";
when 326 => instruction_out <= x"20008200";   -- 0518  IADD32 R0, R1, R0;
when 327 => instruction_out <= x"20008800";   -- 051c  IADD32 R0, R4, R0;
when 328 => instruction_out <= x"30020001";   -- 0520  SHL R0, R0, 0x2; 
when 329 => instruction_out <= x"c4100780";
when 330 => instruction_out <= x"2000c801";   -- 0528  IADD R0, g [0x4], R0; 
when 331 => instruction_out <= x"04200780";
when 332 => instruction_out <= x"d00e0029";   -- 0530  GST.U32 global14[R0], R10; 
when 333 => instruction_out <= x"a0c00781";
when 334 => instruction_out <= x"30000003";   -- RET
when 335 => instruction_out <= x"00000780";

			when others => null;
		end case;
	end process;

end arch;
