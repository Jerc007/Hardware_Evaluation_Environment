

module fence_registers_1_0 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16, n15
;

  DFFR_X1 fence_en_out_reg ( .D(n16), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n10) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n14), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n9) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n13), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n8) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n12), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n7) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n11), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n6) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n1) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n2) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n3) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n4) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n5) );
  OAI21_X1 U2 ( .B1(n6), .B2(cta_id_ld), .A(n1), .ZN(n11) );
  OAI21_X1 U4 ( .B1(n7), .B2(cta_id_ld), .A(n2), .ZN(n12) );
  OAI21_X1 U6 ( .B1(n8), .B2(cta_id_ld), .A(n3), .ZN(n13) );
  OAI21_X1 U8 ( .B1(n9), .B2(cta_id_ld), .A(n4), .ZN(n14) );
  OAI21_X1 U10 ( .B1(n10), .B2(fence_en_ld), .A(n5), .ZN(n16) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_31 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_30 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_29 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_28 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  OAI21_X1 U4 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U6 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U8 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U10 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_27 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_26 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_25 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  OAI21_X1 U4 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U6 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U8 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U10 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_24 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_23 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  OAI21_X1 U4 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U6 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U8 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U10 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_22 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_21 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_20 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_19 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_18 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_17 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_16 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_15 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_14 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_13 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_12 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_11 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_10 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_9 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_8 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_7 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_6 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_5 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_4 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_3 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_2 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  OAI21_X1 U4 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U6 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U8 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U10 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule


module fence_registers_1_1 ( clk_in, host_reset, cta_id_in, cta_id_ld, 
        fence_en_in, fence_en_ld, cta_id_out, fence_en_out );
  input [3:0] cta_id_in;
  output [3:0] cta_id_out;
  input clk_in, host_reset, cta_id_ld, fence_en_in, fence_en_ld;
  output fence_en_out;
  wire   n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31;

  DFFR_X1 fence_en_out_reg ( .D(n17), .CK(clk_in), .RN(n15), .Q(fence_en_out), 
        .QN(n22) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n18), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[3]), .QN(n23) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n19), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[2]), .QN(n24) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n20), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[1]), .QN(n25) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n21), .CK(clk_in), .RN(n15), .Q(
        cta_id_out[0]), .QN(n26) );
  NAND2_X1 U3 ( .A1(cta_id_ld), .A2(cta_id_in[0]), .ZN(n31) );
  NAND2_X1 U5 ( .A1(cta_id_in[1]), .A2(cta_id_ld), .ZN(n30) );
  NAND2_X1 U7 ( .A1(cta_id_in[2]), .A2(cta_id_ld), .ZN(n29) );
  NAND2_X1 U9 ( .A1(cta_id_in[3]), .A2(cta_id_ld), .ZN(n28) );
  NAND2_X1 U12 ( .A1(fence_en_ld), .A2(fence_en_in), .ZN(n27) );
  OAI21_X1 U2 ( .B1(n26), .B2(cta_id_ld), .A(n31), .ZN(n21) );
  OAI21_X1 U4 ( .B1(n25), .B2(cta_id_ld), .A(n30), .ZN(n20) );
  OAI21_X1 U6 ( .B1(n24), .B2(cta_id_ld), .A(n29), .ZN(n19) );
  OAI21_X1 U8 ( .B1(n23), .B2(cta_id_ld), .A(n28), .ZN(n18) );
  OAI21_X1 U10 ( .B1(n22), .B2(fence_en_ld), .A(n27), .ZN(n17) );
  INV_X1 U11 ( .A(host_reset), .ZN(n15) );
endmodule





module warp_checker_SHMEM_ADDR_SIZE14_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, 
        GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  INV_X1 U1 ( .A(A[0]), .ZN(n3) );
  INV_X1 U2 ( .A(A[1]), .ZN(n2) );
  INV_X1 U3 ( .A(B[1]), .ZN(n1) );
  NOR4_X1 U4 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(EQ) );
  NAND4_X1 U5 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .ZN(n7) );
  XNOR2_X1 U6 ( .A(B[3]), .B(A[3]), .ZN(n11) );
  XNOR2_X1 U7 ( .A(B[4]), .B(A[4]), .ZN(n10) );
  XNOR2_X1 U8 ( .A(B[5]), .B(A[5]), .ZN(n9) );
  XNOR2_X1 U9 ( .A(B[6]), .B(A[6]), .ZN(n8) );
  NAND4_X1 U10 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .ZN(n6) );
  OAI22_X1 U11 ( .A1(n16), .A2(n2), .B1(B[1]), .B2(n16), .ZN(n15) );
  AND2_X1 U12 ( .A1(B[0]), .A2(n3), .ZN(n16) );
  OAI22_X1 U13 ( .A1(A[1]), .A2(n17), .B1(n17), .B2(n1), .ZN(n14) );
  NOR2_X1 U14 ( .A1(n3), .A2(B[0]), .ZN(n17) );
  XNOR2_X1 U15 ( .A(B[31]), .B(A[31]), .ZN(n13) );
  XNOR2_X1 U16 ( .A(B[2]), .B(A[2]), .ZN(n12) );
  NAND2_X1 U17 ( .A1(n18), .A2(n19), .ZN(n5) );
  NOR4_X1 U18 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n19) );
  XOR2_X1 U19 ( .A(B[10]), .B(A[10]), .Z(n23) );
  XOR2_X1 U20 ( .A(B[9]), .B(A[9]), .Z(n22) );
  XOR2_X1 U21 ( .A(B[8]), .B(A[8]), .Z(n21) );
  XOR2_X1 U22 ( .A(B[7]), .B(A[7]), .Z(n20) );
  NOR4_X1 U23 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n18) );
  XOR2_X1 U24 ( .A(B[14]), .B(A[14]), .Z(n27) );
  XOR2_X1 U25 ( .A(B[13]), .B(A[13]), .Z(n26) );
  XOR2_X1 U26 ( .A(B[12]), .B(A[12]), .Z(n25) );
  XOR2_X1 U27 ( .A(B[11]), .B(A[11]), .Z(n24) );
  NAND4_X1 U28 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n4) );
  NOR4_X1 U29 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(n31) );
  XOR2_X1 U30 ( .A(B[18]), .B(A[18]), .Z(n35) );
  XOR2_X1 U31 ( .A(B[17]), .B(A[17]), .Z(n34) );
  XOR2_X1 U32 ( .A(B[16]), .B(A[16]), .Z(n33) );
  XOR2_X1 U33 ( .A(B[15]), .B(A[15]), .Z(n32) );
  NOR4_X1 U34 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n30) );
  XOR2_X1 U35 ( .A(B[22]), .B(A[22]), .Z(n39) );
  XOR2_X1 U36 ( .A(B[21]), .B(A[21]), .Z(n38) );
  XOR2_X1 U37 ( .A(B[20]), .B(A[20]), .Z(n37) );
  XOR2_X1 U38 ( .A(B[19]), .B(A[19]), .Z(n36) );
  NOR4_X1 U39 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n29) );
  XOR2_X1 U40 ( .A(B[26]), .B(A[26]), .Z(n43) );
  XOR2_X1 U41 ( .A(B[25]), .B(A[25]), .Z(n42) );
  XOR2_X1 U42 ( .A(B[24]), .B(A[24]), .Z(n41) );
  XOR2_X1 U43 ( .A(B[23]), .B(A[23]), .Z(n40) );
  NOR4_X1 U44 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n28) );
  XOR2_X1 U45 ( .A(B[30]), .B(A[30]), .Z(n47) );
  XOR2_X1 U46 ( .A(B[29]), .B(A[29]), .Z(n46) );
  XOR2_X1 U47 ( .A(B[28]), .B(A[28]), .Z(n45) );
  XOR2_X1 U48 ( .A(B[27]), .B(A[27]), .Z(n44) );
endmodule


module warp_checker ( clk_in, host_reset, reset, en, 
        warp_id_in, warp_lane_id_in, cta_id_in, initial_mask_in, 
        current_mask_in, shmem_base_addr_in, gprs_base_addr_in, next_pc_in, 
        warp_state_in, warps_per_block_in, warp_pool_addr_out, 
        warp_pool_wr_en_out, warp_pool_wr_data_out, warp_state_addr_out, 
        warp_state_wr_en_out, warp_state_wr_data_out, fence_regs_fence_en_out, 
        fence_regs_fence_en_ld, .fence_regs_cta_id_in({
        \fence_regs_cta_id_in[31><3] , \fence_regs_cta_id_in[31><2] , 
        \fence_regs_cta_id_in[31><1] , \fence_regs_cta_id_in[31><0] , 
        \fence_regs_cta_id_in[30><3] , \fence_regs_cta_id_in[30><2] , 
        \fence_regs_cta_id_in[30><1] , \fence_regs_cta_id_in[30><0] , 
        \fence_regs_cta_id_in[29><3] , \fence_regs_cta_id_in[29><2] , 
        \fence_regs_cta_id_in[29><1] , \fence_regs_cta_id_in[29><0] , 
        \fence_regs_cta_id_in[28><3] , \fence_regs_cta_id_in[28><2] , 
        \fence_regs_cta_id_in[28><1] , \fence_regs_cta_id_in[28><0] , 
        \fence_regs_cta_id_in[27><3] , \fence_regs_cta_id_in[27><2] , 
        \fence_regs_cta_id_in[27><1] , \fence_regs_cta_id_in[27><0] , 
        \fence_regs_cta_id_in[26><3] , \fence_regs_cta_id_in[26><2] , 
        \fence_regs_cta_id_in[26><1] , \fence_regs_cta_id_in[26><0] , 
        \fence_regs_cta_id_in[25><3] , \fence_regs_cta_id_in[25><2] , 
        \fence_regs_cta_id_in[25><1] , \fence_regs_cta_id_in[25><0] , 
        \fence_regs_cta_id_in[24><3] , \fence_regs_cta_id_in[24><2] , 
        \fence_regs_cta_id_in[24><1] , \fence_regs_cta_id_in[24><0] , 
        \fence_regs_cta_id_in[23><3] , \fence_regs_cta_id_in[23><2] , 
        \fence_regs_cta_id_in[23><1] , \fence_regs_cta_id_in[23><0] , 
        \fence_regs_cta_id_in[22><3] , \fence_regs_cta_id_in[22><2] , 
        \fence_regs_cta_id_in[22><1] , \fence_regs_cta_id_in[22><0] , 
        \fence_regs_cta_id_in[21><3] , \fence_regs_cta_id_in[21><2] , 
        \fence_regs_cta_id_in[21><1] , \fence_regs_cta_id_in[21><0] , 
        \fence_regs_cta_id_in[20><3] , \fence_regs_cta_id_in[20><2] , 
        \fence_regs_cta_id_in[20><1] , \fence_regs_cta_id_in[20><0] , 
        \fence_regs_cta_id_in[19><3] , \fence_regs_cta_id_in[19><2] , 
        \fence_regs_cta_id_in[19><1] , \fence_regs_cta_id_in[19><0] , 
        \fence_regs_cta_id_in[18><3] , \fence_regs_cta_id_in[18><2] , 
        \fence_regs_cta_id_in[18><1] , \fence_regs_cta_id_in[18><0] , 
        \fence_regs_cta_id_in[17><3] , \fence_regs_cta_id_in[17><2] , 
        \fence_regs_cta_id_in[17><1] , \fence_regs_cta_id_in[17><0] , 
        \fence_regs_cta_id_in[16><3] , \fence_regs_cta_id_in[16><2] , 
        \fence_regs_cta_id_in[16><1] , \fence_regs_cta_id_in[16><0] , 
        \fence_regs_cta_id_in[15><3] , \fence_regs_cta_id_in[15><2] , 
        \fence_regs_cta_id_in[15><1] , \fence_regs_cta_id_in[15><0] , 
        \fence_regs_cta_id_in[14><3] , \fence_regs_cta_id_in[14><2] , 
        \fence_regs_cta_id_in[14><1] , \fence_regs_cta_id_in[14><0] , 
        \fence_regs_cta_id_in[13><3] , \fence_regs_cta_id_in[13><2] , 
        \fence_regs_cta_id_in[13><1] , \fence_regs_cta_id_in[13><0] , 
        \fence_regs_cta_id_in[12><3] , \fence_regs_cta_id_in[12><2] , 
        \fence_regs_cta_id_in[12><1] , \fence_regs_cta_id_in[12><0] , 
        \fence_regs_cta_id_in[11><3] , \fence_regs_cta_id_in[11><2] , 
        \fence_regs_cta_id_in[11><1] , \fence_regs_cta_id_in[11><0] , 
        \fence_regs_cta_id_in[10><3] , \fence_regs_cta_id_in[10><2] , 
        \fence_regs_cta_id_in[10><1] , \fence_regs_cta_id_in[10><0] , 
        \fence_regs_cta_id_in[9><3] , \fence_regs_cta_id_in[9><2] , 
        \fence_regs_cta_id_in[9><1] , \fence_regs_cta_id_in[9><0] , 
        \fence_regs_cta_id_in[8><3] , \fence_regs_cta_id_in[8><2] , 
        \fence_regs_cta_id_in[8><1] , \fence_regs_cta_id_in[8><0] , 
        \fence_regs_cta_id_in[7><3] , \fence_regs_cta_id_in[7><2] , 
        \fence_regs_cta_id_in[7><1] , \fence_regs_cta_id_in[7><0] , 
        \fence_regs_cta_id_in[6><3] , \fence_regs_cta_id_in[6><2] , 
        \fence_regs_cta_id_in[6><1] , \fence_regs_cta_id_in[6><0] , 
        \fence_regs_cta_id_in[5><3] , \fence_regs_cta_id_in[5><2] , 
        \fence_regs_cta_id_in[5><1] , \fence_regs_cta_id_in[5><0] , 
        \fence_regs_cta_id_in[4><3] , \fence_regs_cta_id_in[4><2] , 
        \fence_regs_cta_id_in[4><1] , \fence_regs_cta_id_in[4><0] , 
        \fence_regs_cta_id_in[3><3] , \fence_regs_cta_id_in[3><2] , 
        \fence_regs_cta_id_in[3><1] , \fence_regs_cta_id_in[3><0] , 
        \fence_regs_cta_id_in[2><3] , \fence_regs_cta_id_in[2><2] , 
        \fence_regs_cta_id_in[2><1] , \fence_regs_cta_id_in[2><0] , 
        \fence_regs_cta_id_in[1><3] , \fence_regs_cta_id_in[1><2] , 
        \fence_regs_cta_id_in[1><1] , \fence_regs_cta_id_in[1><0] , 
        \fence_regs_cta_id_in[0><3] , \fence_regs_cta_id_in[0><2] , 
        \fence_regs_cta_id_in[0><1] , \fence_regs_cta_id_in[0><0] }), 
        fence_regs_fence_en_in, warps_done_mask_out, pipeline_stall_out );
  input [4:0] warp_id_in;
  input [1:0] warp_lane_id_in;
  input [3:0] cta_id_in;
  input [31:0] initial_mask_in;
  input [31:0] current_mask_in;
  input [13:0] shmem_base_addr_in;
  input [8:0] gprs_base_addr_in;
  input [31:0] next_pc_in;
  input [1:0] warp_state_in;
  input [5:0] warps_per_block_in;
  output [4:0] warp_pool_addr_out;
  output [127:0] warp_pool_wr_data_out;
  output [4:0] warp_state_addr_out;
  output [1:0] warp_state_wr_data_out;
  output [31:0] fence_regs_fence_en_out;
  output [31:0] fence_regs_fence_en_ld;
  input [31:0] fence_regs_fence_en_in;
  output [31:0] warps_done_mask_out;
  input clk_in, host_reset, reset, en, \fence_regs_cta_id_in[31><3] ,
         \fence_regs_cta_id_in[31><2] , \fence_regs_cta_id_in[31><1] ,
         \fence_regs_cta_id_in[31><0] , \fence_regs_cta_id_in[30><3] ,
         \fence_regs_cta_id_in[30><2] , \fence_regs_cta_id_in[30><1] ,
         \fence_regs_cta_id_in[30><0] , \fence_regs_cta_id_in[29><3] ,
         \fence_regs_cta_id_in[29><2] , \fence_regs_cta_id_in[29><1] ,
         \fence_regs_cta_id_in[29><0] , \fence_regs_cta_id_in[28><3] ,
         \fence_regs_cta_id_in[28><2] , \fence_regs_cta_id_in[28><1] ,
         \fence_regs_cta_id_in[28><0] , \fence_regs_cta_id_in[27><3] ,
         \fence_regs_cta_id_in[27><2] , \fence_regs_cta_id_in[27><1] ,
         \fence_regs_cta_id_in[27><0] , \fence_regs_cta_id_in[26><3] ,
         \fence_regs_cta_id_in[26><2] , \fence_regs_cta_id_in[26><1] ,
         \fence_regs_cta_id_in[26><0] , \fence_regs_cta_id_in[25><3] ,
         \fence_regs_cta_id_in[25><2] , \fence_regs_cta_id_in[25><1] ,
         \fence_regs_cta_id_in[25><0] , \fence_regs_cta_id_in[24><3] ,
         \fence_regs_cta_id_in[24><2] , \fence_regs_cta_id_in[24><1] ,
         \fence_regs_cta_id_in[24><0] , \fence_regs_cta_id_in[23><3] ,
         \fence_regs_cta_id_in[23><2] , \fence_regs_cta_id_in[23><1] ,
         \fence_regs_cta_id_in[23><0] , \fence_regs_cta_id_in[22><3] ,
         \fence_regs_cta_id_in[22><2] , \fence_regs_cta_id_in[22><1] ,
         \fence_regs_cta_id_in[22><0] , \fence_regs_cta_id_in[21><3] ,
         \fence_regs_cta_id_in[21><2] , \fence_regs_cta_id_in[21><1] ,
         \fence_regs_cta_id_in[21><0] , \fence_regs_cta_id_in[20><3] ,
         \fence_regs_cta_id_in[20><2] , \fence_regs_cta_id_in[20><1] ,
         \fence_regs_cta_id_in[20><0] , \fence_regs_cta_id_in[19><3] ,
         \fence_regs_cta_id_in[19><2] , \fence_regs_cta_id_in[19><1] ,
         \fence_regs_cta_id_in[19><0] , \fence_regs_cta_id_in[18><3] ,
         \fence_regs_cta_id_in[18><2] , \fence_regs_cta_id_in[18><1] ,
         \fence_regs_cta_id_in[18><0] , \fence_regs_cta_id_in[17><3] ,
         \fence_regs_cta_id_in[17><2] , \fence_regs_cta_id_in[17><1] ,
         \fence_regs_cta_id_in[17><0] , \fence_regs_cta_id_in[16><3] ,
         \fence_regs_cta_id_in[16><2] , \fence_regs_cta_id_in[16><1] ,
         \fence_regs_cta_id_in[16><0] , \fence_regs_cta_id_in[15><3] ,
         \fence_regs_cta_id_in[15><2] , \fence_regs_cta_id_in[15><1] ,
         \fence_regs_cta_id_in[15><0] , \fence_regs_cta_id_in[14><3] ,
         \fence_regs_cta_id_in[14><2] , \fence_regs_cta_id_in[14><1] ,
         \fence_regs_cta_id_in[14><0] , \fence_regs_cta_id_in[13><3] ,
         \fence_regs_cta_id_in[13><2] , \fence_regs_cta_id_in[13><1] ,
         \fence_regs_cta_id_in[13><0] , \fence_regs_cta_id_in[12><3] ,
         \fence_regs_cta_id_in[12><2] , \fence_regs_cta_id_in[12><1] ,
         \fence_regs_cta_id_in[12><0] , \fence_regs_cta_id_in[11><3] ,
         \fence_regs_cta_id_in[11><2] , \fence_regs_cta_id_in[11><1] ,
         \fence_regs_cta_id_in[11><0] , \fence_regs_cta_id_in[10><3] ,
         \fence_regs_cta_id_in[10><2] , \fence_regs_cta_id_in[10><1] ,
         \fence_regs_cta_id_in[10><0] , \fence_regs_cta_id_in[9><3] ,
         \fence_regs_cta_id_in[9><2] , \fence_regs_cta_id_in[9><1] ,
         \fence_regs_cta_id_in[9><0] , \fence_regs_cta_id_in[8><3] ,
         \fence_regs_cta_id_in[8><2] , \fence_regs_cta_id_in[8><1] ,
         \fence_regs_cta_id_in[8><0] , \fence_regs_cta_id_in[7><3] ,
         \fence_regs_cta_id_in[7><2] , \fence_regs_cta_id_in[7><1] ,
         \fence_regs_cta_id_in[7><0] , \fence_regs_cta_id_in[6><3] ,
         \fence_regs_cta_id_in[6><2] , \fence_regs_cta_id_in[6><1] ,
         \fence_regs_cta_id_in[6><0] , \fence_regs_cta_id_in[5><3] ,
         \fence_regs_cta_id_in[5><2] , \fence_regs_cta_id_in[5><1] ,
         \fence_regs_cta_id_in[5><0] , \fence_regs_cta_id_in[4><3] ,
         \fence_regs_cta_id_in[4><2] , \fence_regs_cta_id_in[4><1] ,
         \fence_regs_cta_id_in[4><0] , \fence_regs_cta_id_in[3><3] ,
         \fence_regs_cta_id_in[3><2] , \fence_regs_cta_id_in[3><1] ,
         \fence_regs_cta_id_in[3><0] , \fence_regs_cta_id_in[2><3] ,
         \fence_regs_cta_id_in[2><2] , \fence_regs_cta_id_in[2><1] ,
         \fence_regs_cta_id_in[2><0] , \fence_regs_cta_id_in[1><3] ,
         \fence_regs_cta_id_in[1><2] , \fence_regs_cta_id_in[1><1] ,
         \fence_regs_cta_id_in[1><0] , \fence_regs_cta_id_in[0><3] ,
         \fence_regs_cta_id_in[0><2] , \fence_regs_cta_id_in[0><1] ,
         \fence_regs_cta_id_in[0><0] ;
  output warp_pool_wr_en_out, warp_state_wr_en_out, pipeline_stall_out;
  wire   N112, N113, N114, N115, N116, \warp_cntr[5] , N567, N572, N703, N704,
         N705, N706, N707, N1190, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         \add_154/carry[5] , \add_154/carry[4] , \add_154/carry[3] ,
         \add_154/carry[2] , n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651;
  wire   [4:0] warp_id_addr;
  wire   [31:0] warps_done_mask;
  wire   [2:0] warp_checker_state_machine;
  wire   [31:0] cta_id_mask_rev;
  wire   [31:0] fence_id_mask;
  assign warp_pool_wr_data_out[127] = 1'b0;
  assign warp_pool_wr_data_out[126] = 1'b0;
  assign warp_pool_wr_data_out[125] = 1'b0;
  assign warp_pool_wr_data_out[124] = 1'b0;
  assign warp_pool_wr_data_out[96] = 1'b0;
  assign N1190 = warps_per_block_in[5];

  DFFR_X1 \warp_checker_state_machine_reg[0]  ( .D(n651), .CK(clk_in), .RN(
        n132), .Q(warp_checker_state_machine[0]), .QN(n3) );
  DFFR_X1 \warp_checker_state_machine_reg[2]  ( .D(n1267), .CK(clk_in), .RN(
        n132), .Q(warp_checker_state_machine[2]), .QN(n8) );
  DFFR_X1 \warp_cntr_reg[5]  ( .D(n983), .CK(clk_in), .RN(n132), .Q(
        \warp_cntr[5] ), .QN(n9) );
  DFFR_X1 \warp_cntr_reg[4]  ( .D(n1261), .CK(clk_in), .RN(n132), .Q(N116), 
        .QN(n985) );
  DFFR_X1 \warp_checker_state_machine_reg[1]  ( .D(n1266), .CK(clk_in), .RN(
        n131), .Q(warp_checker_state_machine[1]), .QN(n7) );
  DFFR_X1 \warp_cntr_reg[3]  ( .D(n1262), .CK(clk_in), .RN(n131), .Q(N115), 
        .QN(n986) );
  DFFR_X1 \warp_cntr_reg[2]  ( .D(n1263), .CK(clk_in), .RN(n131), .Q(N114), 
        .QN(n987) );
  DFFR_X1 \warp_cntr_reg[0]  ( .D(n1264), .CK(clk_in), .RN(n131), .Q(N112), 
        .QN(n989) );
  DFFR_X1 \warp_cntr_reg[1]  ( .D(n1265), .CK(clk_in), .RN(n131), .Q(N113), 
        .QN(n988) );
  DFFR_X1 \warps_done_mask_reg[31]  ( .D(n981), .CK(clk_in), .RN(n131), .Q(
        warps_done_mask[31]), .QN(n10) );
  DFFR_X1 \warps_done_mask_reg[30]  ( .D(n980), .CK(clk_in), .RN(n131), .Q(
        warps_done_mask[30]), .QN(n11) );
  DFFR_X1 \warps_done_mask_reg[29]  ( .D(n979), .CK(clk_in), .RN(n131), .Q(
        warps_done_mask[29]), .QN(n12) );
  DFFR_X1 \warps_done_mask_reg[28]  ( .D(n978), .CK(clk_in), .RN(n131), .Q(
        warps_done_mask[28]), .QN(n13) );
  DFFR_X1 \warps_done_mask_reg[27]  ( .D(n977), .CK(clk_in), .RN(n131), .Q(
        warps_done_mask[27]), .QN(n14) );
  DFFR_X1 \warps_done_mask_reg[26]  ( .D(n976), .CK(clk_in), .RN(n131), .Q(
        warps_done_mask[26]), .QN(n15) );
  DFFR_X1 \warps_done_mask_reg[25]  ( .D(n975), .CK(clk_in), .RN(n131), .Q(
        warps_done_mask[25]), .QN(n16) );
  DFFR_X1 \warps_done_mask_reg[24]  ( .D(n974), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[24]), .QN(n17) );
  DFFR_X1 \warps_done_mask_reg[23]  ( .D(n973), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[23]), .QN(n18) );
  DFFR_X1 \warps_done_mask_reg[22]  ( .D(n972), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[22]), .QN(n19) );
  DFFR_X1 \warps_done_mask_reg[21]  ( .D(n971), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[21]), .QN(n20) );
  DFFR_X1 \warps_done_mask_reg[20]  ( .D(n970), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[20]), .QN(n21) );
  DFFR_X1 \warps_done_mask_reg[19]  ( .D(n969), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[19]), .QN(n22) );
  DFFR_X1 \warps_done_mask_reg[18]  ( .D(n968), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[18]), .QN(n23) );
  DFFR_X1 \warps_done_mask_reg[17]  ( .D(n967), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[17]), .QN(n24) );
  DFFR_X1 \warps_done_mask_reg[16]  ( .D(n966), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[16]), .QN(n25) );
  DFFR_X1 \warps_done_mask_reg[15]  ( .D(n965), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[15]), .QN(n26) );
  DFFR_X1 \warps_done_mask_reg[14]  ( .D(n964), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[14]), .QN(n27) );
  DFFR_X1 \warps_done_mask_reg[13]  ( .D(n963), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[13]), .QN(n28) );
  DFFR_X1 \warps_done_mask_reg[12]  ( .D(n962), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[12]), .QN(n29) );
  DFFR_X1 \warps_done_mask_reg[11]  ( .D(n961), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[11]), .QN(n30) );
  DFFR_X1 \warps_done_mask_reg[10]  ( .D(n960), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[10]), .QN(n31) );
  DFFR_X1 \warps_done_mask_reg[9]  ( .D(n959), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[9]), .QN(n32) );
  DFFR_X1 \warps_done_mask_reg[8]  ( .D(n958), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[8]), .QN(n33) );
  DFFR_X1 \warps_done_mask_reg[7]  ( .D(n957), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[7]), .QN(n34) );
  DFFR_X1 \warps_done_mask_reg[6]  ( .D(n956), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[6]), .QN(n35) );
  DFFR_X1 \warps_done_mask_reg[5]  ( .D(n955), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[5]), .QN(n36) );
  DFFR_X1 \warps_done_mask_reg[4]  ( .D(n954), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[4]), .QN(n37) );
  DFFR_X1 \warps_done_mask_reg[3]  ( .D(n953), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[3]), .QN(n38) );
  DFFR_X1 \warps_done_mask_reg[2]  ( .D(n952), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[2]), .QN(n39) );
  DFFR_X1 \warps_done_mask_reg[1]  ( .D(n951), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[1]), .QN(n40) );
  DFFR_X1 \warps_done_mask_reg[0]  ( .D(n950), .CK(clk_in), .RN(n128), .Q(
        warps_done_mask[0]), .QN(n41) );
  DFFR_X1 \fence_regs_fence_en_out_reg[16]  ( .D(n1189), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[16]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[17]  ( .D(n1190), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[17]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[18]  ( .D(n1191), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[18]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[19]  ( .D(n1192), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[19]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[20]  ( .D(n1193), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[20]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[21]  ( .D(n1194), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[21]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[22]  ( .D(n1195), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[22]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[23]  ( .D(n1196), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[23]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[24]  ( .D(n1197), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[24]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[25]  ( .D(n1198), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[25]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[26]  ( .D(n1199), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[26]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[27]  ( .D(n1200), .CK(clk_in), .RN(n127), .Q(fence_regs_fence_en_out[27]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[28]  ( .D(n1201), .CK(clk_in), .RN(n127), .Q(fence_regs_fence_en_out[28]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[29]  ( .D(n1202), .CK(clk_in), .RN(n127), .Q(fence_regs_fence_en_out[29]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[30]  ( .D(n1203), .CK(clk_in), .RN(n127), .Q(fence_regs_fence_en_out[30]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[31]  ( .D(n1204), .CK(clk_in), .RN(n127), .Q(fence_regs_fence_en_out[31]) );
  DFFR_X1 \warp_id_addr_reg[1]  ( .D(n1256), .CK(clk_in), .RN(n127), .Q(
        warp_id_addr[1]), .QN(n5) );
  DFFR_X1 \warp_id_addr_reg[2]  ( .D(n1257), .CK(clk_in), .RN(n127), .Q(
        warp_id_addr[2]) );
  DFFR_X1 \warp_id_addr_reg[3]  ( .D(n1258), .CK(clk_in), .RN(n127), .Q(
        warp_id_addr[3]), .QN(n6) );
  DFFR_X1 \warp_id_addr_reg[4]  ( .D(n1259), .CK(clk_in), .RN(n127), .Q(
        warp_id_addr[4]) );
  DFFR_X1 \warp_id_addr_reg[0]  ( .D(n1260), .CK(clk_in), .RN(n127), .Q(
        warp_id_addr[0]), .QN(n4) );
  DFFR_X1 pipeline_stall_out_reg ( .D(n1255), .CK(clk_in), .RN(n127), .Q(
        pipeline_stall_out) );
  DFFR_X1 \warps_done_mask_out_reg[31]  ( .D(n1109), .CK(clk_in), .RN(n127), 
        .Q(warps_done_mask_out[31]) );
  DFFR_X1 \warps_done_mask_out_reg[30]  ( .D(n1110), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[30]) );
  DFFR_X1 \warps_done_mask_out_reg[29]  ( .D(n1111), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[29]) );
  DFFR_X1 \warps_done_mask_out_reg[28]  ( .D(n1112), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[28]) );
  DFFR_X1 \warps_done_mask_out_reg[27]  ( .D(n1113), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[27]) );
  DFFR_X1 \warps_done_mask_out_reg[26]  ( .D(n1114), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[26]) );
  DFFR_X1 \warps_done_mask_out_reg[25]  ( .D(n1115), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[25]) );
  DFFR_X1 \warps_done_mask_out_reg[24]  ( .D(n1116), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[24]) );
  DFFR_X1 \warps_done_mask_out_reg[23]  ( .D(n1117), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[23]) );
  DFFR_X1 \warps_done_mask_out_reg[22]  ( .D(n1118), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[22]) );
  DFFR_X1 \warps_done_mask_out_reg[21]  ( .D(n1119), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[21]) );
  DFFR_X1 \warps_done_mask_out_reg[20]  ( .D(n1120), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[20]) );
  DFFR_X1 \warps_done_mask_out_reg[19]  ( .D(n1121), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[19]) );
  DFFR_X1 \warps_done_mask_out_reg[18]  ( .D(n1122), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[18]) );
  DFFR_X1 \warps_done_mask_out_reg[17]  ( .D(n1123), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[17]) );
  DFFR_X1 \warps_done_mask_out_reg[16]  ( .D(n1124), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[16]) );
  DFFR_X1 \warps_done_mask_out_reg[15]  ( .D(n1125), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[15]) );
  DFFR_X1 \warps_done_mask_out_reg[14]  ( .D(n1126), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[14]) );
  DFFR_X1 \warps_done_mask_out_reg[13]  ( .D(n1127), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[13]) );
  DFFR_X1 \warps_done_mask_out_reg[12]  ( .D(n1128), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[12]) );
  DFFR_X1 \warps_done_mask_out_reg[11]  ( .D(n1129), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[11]) );
  DFFR_X1 \warps_done_mask_out_reg[10]  ( .D(n1130), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[10]) );
  DFFR_X1 \warps_done_mask_out_reg[9]  ( .D(n1131), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[9]) );
  DFFR_X1 \warps_done_mask_out_reg[8]  ( .D(n1132), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[8]) );
  DFFR_X1 \warps_done_mask_out_reg[7]  ( .D(n1133), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[7]) );
  DFFR_X1 \warps_done_mask_out_reg[6]  ( .D(n1134), .CK(clk_in), .RN(n124), 
        .Q(warps_done_mask_out[6]) );
  DFFR_X1 \warps_done_mask_out_reg[5]  ( .D(n1135), .CK(clk_in), .RN(n124), 
        .Q(warps_done_mask_out[5]) );
  DFFR_X1 \warps_done_mask_out_reg[4]  ( .D(n1136), .CK(clk_in), .RN(n124), 
        .Q(warps_done_mask_out[4]) );
  DFFR_X1 \warps_done_mask_out_reg[3]  ( .D(n1137), .CK(clk_in), .RN(n124), 
        .Q(warps_done_mask_out[3]) );
  DFFR_X1 \warps_done_mask_out_reg[2]  ( .D(n1138), .CK(clk_in), .RN(n124), 
        .Q(warps_done_mask_out[2]) );
  DFFR_X1 \warps_done_mask_out_reg[1]  ( .D(n1139), .CK(clk_in), .RN(n124), 
        .Q(warps_done_mask_out[1]) );
  DFFR_X1 \warps_done_mask_out_reg[0]  ( .D(n1140), .CK(clk_in), .RN(n124), 
        .Q(warps_done_mask_out[0]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[23]  ( .D(n1231), .CK(clk_in), .RN(n124), 
        .Q(fence_regs_fence_en_ld[23]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[22]  ( .D(n1232), .CK(clk_in), .RN(n124), 
        .Q(fence_regs_fence_en_ld[22]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[21]  ( .D(n1233), .CK(clk_in), .RN(n124), 
        .Q(fence_regs_fence_en_ld[21]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[20]  ( .D(n1234), .CK(clk_in), .RN(n124), 
        .Q(fence_regs_fence_en_ld[20]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[19]  ( .D(n1235), .CK(clk_in), .RN(n124), 
        .Q(fence_regs_fence_en_ld[19]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[18]  ( .D(n1236), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[18]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[17]  ( .D(n1237), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[17]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[16]  ( .D(n1238), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[16]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[31]  ( .D(n1223), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[31]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[30]  ( .D(n1224), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[30]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[29]  ( .D(n1225), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[29]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[28]  ( .D(n1226), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[28]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[27]  ( .D(n1227), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[27]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[26]  ( .D(n1228), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[26]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[25]  ( .D(n1229), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[25]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[24]  ( .D(n1230), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[24]) );
  DFFR_X1 warp_pool_wr_en_out_reg ( .D(n1216), .CK(clk_in), .RN(n123), .Q(
        warp_pool_wr_en_out), .QN(n787) );
  DFFR_X1 \warp_pool_addr_out_reg[2]  ( .D(n1213), .CK(clk_in), .RN(n122), .Q(
        warp_pool_addr_out[2]), .QN(n790) );
  DFFR_X1 \warp_pool_addr_out_reg[3]  ( .D(n1214), .CK(clk_in), .RN(n122), .Q(
        warp_pool_addr_out[3]), .QN(n789) );
  DFFR_X1 \warp_pool_addr_out_reg[4]  ( .D(n1215), .CK(clk_in), .RN(n122), .Q(
        warp_pool_addr_out[4]), .QN(n788) );
  DFFR_X1 \warp_pool_addr_out_reg[1]  ( .D(n1217), .CK(clk_in), .RN(n122), .Q(
        warp_pool_addr_out[1]), .QN(n786) );
  DFFR_X1 \warp_pool_wr_data_out_reg[106]  ( .D(n1218), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[106]), .QN(n785) );
  DFFR_X1 \warp_pool_wr_data_out_reg[107]  ( .D(n1219), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[107]), .QN(n784) );
  DFFR_X1 \warp_pool_wr_data_out_reg[108]  ( .D(n1220), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[108]), .QN(n783) );
  DFFR_X1 \warp_pool_wr_data_out_reg[109]  ( .D(n1221), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[109]), .QN(n782) );
  DFFR_X1 \warp_pool_addr_out_reg[0]  ( .D(n1222), .CK(clk_in), .RN(n122), .Q(
        warp_pool_addr_out[0]), .QN(n781) );
  DFFR_X1 warp_state_wr_en_out_reg ( .D(n1206), .CK(clk_in), .RN(n122), .Q(
        warp_state_wr_en_out), .QN(n796) );
  DFFR_X1 \warp_state_addr_out_reg[1]  ( .D(n1207), .CK(clk_in), .RN(n122), 
        .Q(warp_state_addr_out[1]), .QN(n795) );
  DFFR_X1 \warp_state_addr_out_reg[2]  ( .D(n1208), .CK(clk_in), .RN(n122), 
        .Q(warp_state_addr_out[2]), .QN(n794) );
  DFFR_X1 \warp_state_addr_out_reg[3]  ( .D(n1209), .CK(clk_in), .RN(n121), 
        .Q(warp_state_addr_out[3]), .QN(n793) );
  DFFR_X1 \warp_state_wr_data_out_reg[0]  ( .D(n1211), .CK(clk_in), .RN(n121), 
        .Q(warp_state_wr_data_out[0]), .QN(n1173) );
  DFFR_X1 \warp_state_addr_out_reg[0]  ( .D(n1212), .CK(clk_in), .RN(n121), 
        .Q(warp_state_addr_out[0]), .QN(n791) );
  DFFR_X1 \warp_state_wr_data_out_reg[1]  ( .D(n984), .CK(clk_in), .RN(n121), 
        .Q(warp_state_wr_data_out[1]), .QN(n917) );
  DFFR_X1 \warp_pool_wr_data_out_reg[0]  ( .D(n1108), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[0]), .QN(n916) );
  DFFR_X1 \warp_pool_wr_data_out_reg[1]  ( .D(n1107), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[1]), .QN(n915) );
  DFFR_X1 \warp_pool_wr_data_out_reg[2]  ( .D(n1106), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[2]), .QN(n914) );
  DFFR_X1 \warp_pool_wr_data_out_reg[3]  ( .D(n1105), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[3]), .QN(n913) );
  DFFR_X1 \warp_pool_wr_data_out_reg[4]  ( .D(n1104), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[4]), .QN(n912) );
  DFFR_X1 \warp_pool_wr_data_out_reg[5]  ( .D(n1103), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[5]), .QN(n911) );
  DFFR_X1 \warp_pool_wr_data_out_reg[6]  ( .D(n1102), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[6]), .QN(n910) );
  DFFR_X1 \warp_pool_wr_data_out_reg[7]  ( .D(n1101), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[7]), .QN(n909) );
  DFFR_X1 \warp_pool_wr_data_out_reg[8]  ( .D(n1100), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[8]), .QN(n908) );
  DFFR_X1 \warp_pool_wr_data_out_reg[9]  ( .D(n1099), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[9]), .QN(n907) );
  DFFR_X1 \warp_pool_wr_data_out_reg[10]  ( .D(n1098), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[10]), .QN(n906) );
  DFFR_X1 \warp_pool_wr_data_out_reg[11]  ( .D(n1097), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[11]), .QN(n905) );
  DFFR_X1 \warp_pool_wr_data_out_reg[12]  ( .D(n1096), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[12]), .QN(n904) );
  DFFR_X1 \warp_pool_wr_data_out_reg[13]  ( .D(n1095), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[13]), .QN(n903) );
  DFFR_X1 \warp_pool_wr_data_out_reg[14]  ( .D(n1094), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[14]), .QN(n902) );
  DFFR_X1 \warp_pool_wr_data_out_reg[15]  ( .D(n1093), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[15]), .QN(n901) );
  DFFR_X1 \warp_pool_wr_data_out_reg[16]  ( .D(n1092), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[16]), .QN(n900) );
  DFFR_X1 \warp_pool_wr_data_out_reg[17]  ( .D(n1091), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[17]), .QN(n899) );
  DFFR_X1 \warp_pool_wr_data_out_reg[18]  ( .D(n1090), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[18]), .QN(n898) );
  DFFR_X1 \warp_pool_wr_data_out_reg[19]  ( .D(n1089), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[19]), .QN(n897) );
  DFFR_X1 \warp_pool_wr_data_out_reg[20]  ( .D(n1088), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[20]), .QN(n896) );
  DFFR_X1 \warp_pool_wr_data_out_reg[21]  ( .D(n1087), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[21]), .QN(n895) );
  DFFR_X1 \warp_pool_wr_data_out_reg[22]  ( .D(n1086), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[22]), .QN(n894) );
  DFFR_X1 \warp_pool_wr_data_out_reg[23]  ( .D(n1085), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[23]), .QN(n893) );
  DFFR_X1 \warp_pool_wr_data_out_reg[24]  ( .D(n1084), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[24]), .QN(n892) );
  DFFR_X1 \warp_pool_wr_data_out_reg[25]  ( .D(n1083), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[25]), .QN(n891) );
  DFFR_X1 \warp_pool_wr_data_out_reg[26]  ( .D(n1082), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[26]), .QN(n890) );
  DFFR_X1 \warp_pool_wr_data_out_reg[27]  ( .D(n1081), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[27]), .QN(n889) );
  DFFR_X1 \warp_pool_wr_data_out_reg[28]  ( .D(n1080), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[28]), .QN(n888) );
  DFFR_X1 \warp_pool_wr_data_out_reg[29]  ( .D(n1079), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[29]), .QN(n887) );
  DFFR_X1 \warp_pool_wr_data_out_reg[30]  ( .D(n1078), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[30]), .QN(n886) );
  DFFR_X1 \warp_pool_wr_data_out_reg[31]  ( .D(n1077), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[31]), .QN(n885) );
  DFFR_X1 \warp_pool_wr_data_out_reg[32]  ( .D(n1076), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[32]), .QN(n884) );
  DFFR_X1 \warp_pool_wr_data_out_reg[33]  ( .D(n1075), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[33]), .QN(n883) );
  DFFR_X1 \warp_pool_wr_data_out_reg[34]  ( .D(n1074), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[34]), .QN(n882) );
  DFFR_X1 \warp_pool_wr_data_out_reg[35]  ( .D(n1073), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[35]), .QN(n881) );
  DFFR_X1 \warp_pool_wr_data_out_reg[36]  ( .D(n1072), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[36]), .QN(n880) );
  DFFR_X1 \warp_pool_wr_data_out_reg[37]  ( .D(n1071), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[37]), .QN(n879) );
  DFFR_X1 \warp_pool_wr_data_out_reg[38]  ( .D(n1070), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[38]), .QN(n878) );
  DFFR_X1 \warp_pool_wr_data_out_reg[39]  ( .D(n1069), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[39]), .QN(n877) );
  DFFR_X1 \warp_pool_wr_data_out_reg[40]  ( .D(n1068), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[40]), .QN(n876) );
  DFFR_X1 \warp_pool_wr_data_out_reg[41]  ( .D(n1067), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[41]), .QN(n875) );
  DFFR_X1 \warp_pool_wr_data_out_reg[42]  ( .D(n1066), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[42]), .QN(n874) );
  DFFR_X1 \warp_pool_wr_data_out_reg[43]  ( .D(n1065), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[43]), .QN(n873) );
  DFFR_X1 \warp_pool_wr_data_out_reg[44]  ( .D(n1064), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[44]), .QN(n872) );
  DFFR_X1 \warp_pool_wr_data_out_reg[45]  ( .D(n1063), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[45]), .QN(n871) );
  DFFR_X1 \warp_pool_wr_data_out_reg[46]  ( .D(n1062), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[46]), .QN(n870) );
  DFFR_X1 \warp_pool_wr_data_out_reg[47]  ( .D(n1061), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[47]), .QN(n869) );
  DFFR_X1 \warp_pool_wr_data_out_reg[48]  ( .D(n1060), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[48]), .QN(n868) );
  DFFR_X1 \warp_pool_wr_data_out_reg[49]  ( .D(n1059), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[49]), .QN(n867) );
  DFFR_X1 \warp_pool_wr_data_out_reg[50]  ( .D(n1058), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[50]), .QN(n866) );
  DFFR_X1 \warp_pool_wr_data_out_reg[51]  ( .D(n1057), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[51]), .QN(n865) );
  DFFR_X1 \warp_pool_wr_data_out_reg[52]  ( .D(n1056), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[52]), .QN(n864) );
  DFFR_X1 \warp_pool_wr_data_out_reg[53]  ( .D(n1055), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[53]), .QN(n863) );
  DFFR_X1 \warp_pool_wr_data_out_reg[54]  ( .D(n1054), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[54]), .QN(n862) );
  DFFR_X1 \warp_pool_wr_data_out_reg[55]  ( .D(n1053), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[55]), .QN(n861) );
  DFFR_X1 \warp_pool_wr_data_out_reg[56]  ( .D(n1052), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[56]), .QN(n860) );
  DFFR_X1 \warp_pool_wr_data_out_reg[57]  ( .D(n1051), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[57]), .QN(n859) );
  DFFR_X1 \warp_pool_wr_data_out_reg[58]  ( .D(n1050), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[58]), .QN(n858) );
  DFFR_X1 \warp_pool_wr_data_out_reg[59]  ( .D(n1049), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[59]), .QN(n857) );
  DFFR_X1 \warp_pool_wr_data_out_reg[60]  ( .D(n1048), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[60]), .QN(n856) );
  DFFR_X1 \warp_pool_wr_data_out_reg[61]  ( .D(n1047), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[61]), .QN(n855) );
  DFFR_X1 \warp_pool_wr_data_out_reg[62]  ( .D(n1046), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[62]), .QN(n854) );
  DFFR_X1 \warp_pool_wr_data_out_reg[63]  ( .D(n1045), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[63]), .QN(n853) );
  DFFR_X1 \warp_pool_wr_data_out_reg[64]  ( .D(n1044), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[64]), .QN(n852) );
  DFFR_X1 \warp_pool_wr_data_out_reg[65]  ( .D(n1043), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[65]), .QN(n851) );
  DFFR_X1 \warp_pool_wr_data_out_reg[66]  ( .D(n1042), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[66]), .QN(n850) );
  DFFR_X1 \warp_pool_wr_data_out_reg[67]  ( .D(n1041), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[67]), .QN(n849) );
  DFFR_X1 \warp_pool_wr_data_out_reg[68]  ( .D(n1040), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[68]), .QN(n848) );
  DFFR_X1 \warp_pool_wr_data_out_reg[69]  ( .D(n1039), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[69]), .QN(n847) );
  DFFR_X1 \warp_pool_wr_data_out_reg[70]  ( .D(n1038), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[70]), .QN(n846) );
  DFFR_X1 \warp_pool_wr_data_out_reg[71]  ( .D(n1037), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[71]), .QN(n845) );
  DFFR_X1 \warp_pool_wr_data_out_reg[72]  ( .D(n1036), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[72]), .QN(n844) );
  DFFR_X1 \warp_pool_wr_data_out_reg[73]  ( .D(n1035), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[73]), .QN(n843) );
  DFFR_X1 \warp_pool_wr_data_out_reg[74]  ( .D(n1034), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[74]), .QN(n842) );
  DFFR_X1 \warp_pool_wr_data_out_reg[75]  ( .D(n1033), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[75]), .QN(n841) );
  DFFR_X1 \warp_pool_wr_data_out_reg[76]  ( .D(n1032), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[76]), .QN(n840) );
  DFFR_X1 \warp_pool_wr_data_out_reg[77]  ( .D(n1031), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[77]), .QN(n839) );
  DFFR_X1 \warp_pool_wr_data_out_reg[78]  ( .D(n1030), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[78]), .QN(n838) );
  DFFR_X1 \warp_pool_wr_data_out_reg[79]  ( .D(n1029), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[79]), .QN(n837) );
  DFFR_X1 \warp_pool_wr_data_out_reg[80]  ( .D(n1028), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[80]), .QN(n836) );
  DFFR_X1 \warp_pool_wr_data_out_reg[81]  ( .D(n1027), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[81]), .QN(n835) );
  DFFR_X1 \warp_pool_wr_data_out_reg[82]  ( .D(n1026), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[82]), .QN(n834) );
  DFFR_X1 \warp_pool_wr_data_out_reg[83]  ( .D(n1025), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[83]), .QN(n833) );
  DFFR_X1 \warp_pool_wr_data_out_reg[84]  ( .D(n1024), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[84]), .QN(n832) );
  DFFR_X1 \warp_pool_wr_data_out_reg[85]  ( .D(n1023), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[85]), .QN(n831) );
  DFFR_X1 \warp_pool_wr_data_out_reg[86]  ( .D(n1022), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[86]), .QN(n830) );
  DFFR_X1 \warp_pool_wr_data_out_reg[87]  ( .D(n1021), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[87]), .QN(n829) );
  DFFR_X1 \warp_pool_wr_data_out_reg[88]  ( .D(n1020), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[88]), .QN(n828) );
  DFFR_X1 \warp_pool_wr_data_out_reg[89]  ( .D(n1019), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[89]), .QN(n827) );
  DFFR_X1 \warp_pool_wr_data_out_reg[90]  ( .D(n1018), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[90]), .QN(n826) );
  DFFR_X1 \warp_pool_wr_data_out_reg[91]  ( .D(n1017), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[91]), .QN(n825) );
  DFFR_X1 \warp_pool_wr_data_out_reg[92]  ( .D(n1016), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[92]), .QN(n824) );
  DFFR_X1 \warp_pool_wr_data_out_reg[93]  ( .D(n1015), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[93]), .QN(n823) );
  DFFR_X1 \warp_pool_wr_data_out_reg[94]  ( .D(n1014), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[94]), .QN(n822) );
  DFFR_X1 \warp_pool_wr_data_out_reg[95]  ( .D(n1013), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[95]), .QN(n821) );
  DFFR_X1 \warp_pool_wr_data_out_reg[97]  ( .D(n1012), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[97]), .QN(n820) );
  DFFR_X1 \warp_pool_wr_data_out_reg[98]  ( .D(n1011), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[98]), .QN(n819) );
  DFFR_X1 \warp_pool_wr_data_out_reg[99]  ( .D(n1010), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[99]), .QN(n818) );
  DFFR_X1 \warp_pool_wr_data_out_reg[100]  ( .D(n1009), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[100]), .QN(n817) );
  DFFR_X1 \warp_pool_wr_data_out_reg[101]  ( .D(n1008), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[101]), .QN(n816) );
  DFFR_X1 \warp_pool_wr_data_out_reg[102]  ( .D(n1007), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[102]), .QN(n815) );
  DFFR_X1 \warp_pool_wr_data_out_reg[103]  ( .D(n1006), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[103]), .QN(n814) );
  DFFR_X1 \warp_pool_wr_data_out_reg[104]  ( .D(n1005), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[104]), .QN(n813) );
  DFFR_X1 \warp_pool_wr_data_out_reg[105]  ( .D(n1004), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[105]), .QN(n812) );
  DFFR_X1 \warp_pool_wr_data_out_reg[110]  ( .D(n1003), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[110]), .QN(n811) );
  DFFR_X1 \warp_pool_wr_data_out_reg[111]  ( .D(n1002), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[111]), .QN(n810) );
  DFFR_X1 \warp_pool_wr_data_out_reg[112]  ( .D(n1001), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[112]), .QN(n809) );
  DFFR_X1 \warp_pool_wr_data_out_reg[113]  ( .D(n1000), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[113]), .QN(n808) );
  DFFR_X1 \warp_pool_wr_data_out_reg[114]  ( .D(n999), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[114]), .QN(n807) );
  DFFR_X1 \warp_pool_wr_data_out_reg[115]  ( .D(n998), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[115]), .QN(n806) );
  DFFR_X1 \warp_pool_wr_data_out_reg[116]  ( .D(n997), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[116]), .QN(n805) );
  DFFR_X1 \warp_pool_wr_data_out_reg[117]  ( .D(n996), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[117]), .QN(n804) );
  DFFR_X1 \warp_pool_wr_data_out_reg[118]  ( .D(n995), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[118]), .QN(n803) );
  DFFR_X1 \warp_pool_wr_data_out_reg[119]  ( .D(n994), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[119]), .QN(n802) );
  DFFR_X1 \warp_pool_wr_data_out_reg[120]  ( .D(n993), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[120]), .QN(n801) );
  DFFR_X1 \warp_pool_wr_data_out_reg[121]  ( .D(n992), .CK(clk_in), .RN(n111), 
        .Q(warp_pool_wr_data_out[121]), .QN(n800) );
  DFFR_X1 \warp_pool_wr_data_out_reg[122]  ( .D(n991), .CK(clk_in), .RN(n111), 
        .Q(warp_pool_wr_data_out[122]), .QN(n799) );
  DFFR_X1 \warp_pool_wr_data_out_reg[123]  ( .D(n990), .CK(clk_in), .RN(n111), 
        .Q(warp_pool_wr_data_out[123]), .QN(n798) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[7]  ( .D(n1247), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_ld[7]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[7]  ( .D(n1180), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_out[7]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[6]  ( .D(n1248), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_ld[6]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[6]  ( .D(n1179), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_out[6]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[5]  ( .D(n1249), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_ld[5]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[5]  ( .D(n1178), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_out[5]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[4]  ( .D(n1250), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_ld[4]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[4]  ( .D(n1177), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_out[4]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[3]  ( .D(n1251), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_ld[3]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[3]  ( .D(n1176), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_out[3]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[2]  ( .D(n1252), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_ld[2]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[2]  ( .D(n1175), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_out[2]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[1]  ( .D(n1253), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_ld[1]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[1]  ( .D(n1174), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_out[1]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[0]  ( .D(n1254), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_ld[0]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[0]  ( .D(n1205), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_out[0]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[15]  ( .D(n1239), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_ld[15]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[15]  ( .D(n1188), .CK(clk_in), .RN(n110), .Q(fence_regs_fence_en_out[15]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[14]  ( .D(n1240), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_ld[14]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[14]  ( .D(n1187), .CK(clk_in), .RN(n110), .Q(fence_regs_fence_en_out[14]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[13]  ( .D(n1241), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_ld[13]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[13]  ( .D(n1186), .CK(clk_in), .RN(n109), .Q(fence_regs_fence_en_out[13]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[12]  ( .D(n1242), .CK(clk_in), .RN(n109), 
        .Q(fence_regs_fence_en_ld[12]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[12]  ( .D(n1185), .CK(clk_in), .RN(n109), .Q(fence_regs_fence_en_out[12]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[11]  ( .D(n1243), .CK(clk_in), .RN(n109), 
        .Q(fence_regs_fence_en_ld[11]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[11]  ( .D(n1184), .CK(clk_in), .RN(n109), .Q(fence_regs_fence_en_out[11]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[10]  ( .D(n1244), .CK(clk_in), .RN(n109), 
        .Q(fence_regs_fence_en_ld[10]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[10]  ( .D(n1183), .CK(clk_in), .RN(n109), .Q(fence_regs_fence_en_out[10]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[9]  ( .D(n1245), .CK(clk_in), .RN(n109), 
        .Q(fence_regs_fence_en_ld[9]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[9]  ( .D(n1182), .CK(clk_in), .RN(n109), 
        .Q(fence_regs_fence_en_out[9]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[8]  ( .D(n1246), .CK(clk_in), .RN(n109), 
        .Q(fence_regs_fence_en_ld[8]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[8]  ( .D(n1181), .CK(clk_in), .RN(n109), 
        .Q(fence_regs_fence_en_out[8]) );
  DFFR_X1 \warp_state_addr_out_reg[4]  ( .D(n1210), .CK(clk_in), .RN(n109), 
        .Q(warp_state_addr_out[4]), .QN(n792) );
  warp_checker_SHMEM_ADDR_SIZE14_DW01_cmp6_0 eq_137 ( .A(cta_id_mask_rev), .B(
        fence_id_mask), .TC(1'b0), .EQ(N567) );
  HA_X1 \add_154/U1_1_1  ( .A(N113), .B(N112), .CO(\add_154/carry[2] ), .S(
        N703) );
  HA_X1 \add_154/U1_1_2  ( .A(N114), .B(\add_154/carry[2] ), .CO(
        \add_154/carry[3] ), .S(N704) );
  HA_X1 \add_154/U1_1_3  ( .A(N115), .B(\add_154/carry[3] ), .CO(
        \add_154/carry[4] ), .S(N705) );
  HA_X1 \add_154/U1_1_4  ( .A(N116), .B(\add_154/carry[4] ), .CO(
        \add_154/carry[5] ), .S(N706) );
  AND3_X1 U3 ( .A1(n197), .A2(n187), .A3(n414), .ZN(n1) );
  NOR3_X2 U4 ( .A1(n6), .A2(warp_id_addr[4]), .A3(n187), .ZN(n224) );
  NOR3_X2 U5 ( .A1(warp_id_addr[3]), .A2(warp_id_addr[4]), .A3(n187), .ZN(n200) );
  BUF_X1 U6 ( .A(n94), .Z(n89) );
  BUF_X1 U7 ( .A(n94), .Z(n88) );
  BUF_X1 U9 ( .A(n94), .Z(n93) );
  BUF_X1 U10 ( .A(n95), .Z(n87) );
  BUF_X1 U11 ( .A(n95), .Z(n86) );
  BUF_X1 U12 ( .A(n95), .Z(n85) );
  BUF_X1 U13 ( .A(n95), .Z(n84) );
  BUF_X1 U14 ( .A(n94), .Z(n92) );
  BUF_X1 U15 ( .A(n94), .Z(n91) );
  BUF_X1 U16 ( .A(n94), .Z(n90) );
  BUF_X1 U17 ( .A(n95), .Z(n83) );
  INV_X1 U18 ( .A(n1), .ZN(n82) );
  INV_X1 U19 ( .A(n1), .ZN(n79) );
  BUF_X1 U20 ( .A(n163), .Z(n96) );
  BUF_X1 U21 ( .A(n163), .Z(n97) );
  BUF_X1 U22 ( .A(n149), .Z(n94) );
  BUF_X1 U23 ( .A(n163), .Z(n98) );
  BUF_X1 U24 ( .A(n149), .Z(n95) );
  BUF_X1 U25 ( .A(n108), .Z(n136) );
  BUF_X1 U26 ( .A(n108), .Z(n135) );
  BUF_X1 U27 ( .A(n107), .Z(n134) );
  BUF_X1 U28 ( .A(n107), .Z(n133) );
  INV_X1 U29 ( .A(n102), .ZN(n100) );
  INV_X1 U30 ( .A(n102), .ZN(n99) );
  BUF_X1 U31 ( .A(n103), .Z(n105) );
  BUF_X1 U32 ( .A(n103), .Z(n104) );
  BUF_X1 U33 ( .A(n103), .Z(n106) );
  BUF_X1 U34 ( .A(n982), .Z(n108) );
  BUF_X1 U35 ( .A(n982), .Z(n107) );
  INV_X1 U36 ( .A(n138), .ZN(n137) );
  INV_X1 U37 ( .A(n140), .ZN(n139) );
  INV_X1 U38 ( .A(n142), .ZN(n141) );
  INV_X1 U39 ( .A(n144), .ZN(n143) );
  INV_X1 U40 ( .A(n53), .ZN(n73) );
  INV_X1 U41 ( .A(n47), .ZN(n71) );
  INV_X1 U42 ( .A(n54), .ZN(n74) );
  NAND2_X1 U43 ( .A1(n1), .A2(n281), .ZN(n160) );
  INV_X1 U44 ( .A(n44), .ZN(n70) );
  INV_X1 U45 ( .A(n60), .ZN(n76) );
  INV_X1 U46 ( .A(n57), .ZN(n75) );
  BUF_X1 U47 ( .A(n42), .Z(n102) );
  BUF_X1 U48 ( .A(n42), .Z(n101) );
  BUF_X1 U49 ( .A(n303), .Z(n103) );
  INV_X1 U50 ( .A(n43), .ZN(n69) );
  INV_X1 U51 ( .A(n48), .ZN(n72) );
  INV_X1 U52 ( .A(cta_id_in[1]), .ZN(n140) );
  INV_X1 U53 ( .A(cta_id_in[3]), .ZN(n144) );
  INV_X1 U54 ( .A(cta_id_in[2]), .ZN(n142) );
  INV_X1 U55 ( .A(cta_id_in[0]), .ZN(n138) );
  OR3_X1 U56 ( .A1(warp_checker_state_machine[1]), .A2(
        warp_checker_state_machine[2]), .A3(warp_checker_state_machine[0]), 
        .ZN(n42) );
  NOR2_X1 U57 ( .A1(n988), .A2(N112), .ZN(n62) );
  NOR2_X1 U58 ( .A1(n988), .A2(n989), .ZN(n61) );
  NOR2_X1 U59 ( .A1(N112), .A2(N113), .ZN(n59) );
  NOR2_X1 U60 ( .A1(n989), .A2(N113), .ZN(n58) );
  AOI22_X1 U61 ( .A1(cta_id_mask_rev[28]), .A2(n59), .B1(cta_id_mask_rev[29]), 
        .B2(n58), .ZN(n43) );
  AOI221_X1 U62 ( .B1(cta_id_mask_rev[30]), .B2(n62), .C1(cta_id_mask_rev[31]), 
        .C2(n61), .A(n69), .ZN(n46) );
  AOI22_X1 U63 ( .A1(cta_id_mask_rev[24]), .A2(n59), .B1(cta_id_mask_rev[25]), 
        .B2(n58), .ZN(n44) );
  AOI221_X1 U64 ( .B1(cta_id_mask_rev[26]), .B2(n62), .C1(cta_id_mask_rev[27]), 
        .C2(n61), .A(n70), .ZN(n45) );
  OAI22_X1 U65 ( .A1(n987), .A2(n46), .B1(N114), .B2(n45), .ZN(n52) );
  AOI22_X1 U66 ( .A1(cta_id_mask_rev[20]), .A2(n59), .B1(cta_id_mask_rev[21]), 
        .B2(n58), .ZN(n47) );
  AOI221_X1 U67 ( .B1(cta_id_mask_rev[22]), .B2(n62), .C1(cta_id_mask_rev[23]), 
        .C2(n61), .A(n71), .ZN(n50) );
  AOI22_X1 U68 ( .A1(cta_id_mask_rev[16]), .A2(n59), .B1(cta_id_mask_rev[17]), 
        .B2(n58), .ZN(n48) );
  AOI221_X1 U69 ( .B1(cta_id_mask_rev[18]), .B2(n62), .C1(cta_id_mask_rev[19]), 
        .C2(n61), .A(n72), .ZN(n49) );
  OAI22_X1 U70 ( .A1(n50), .A2(n987), .B1(N114), .B2(n49), .ZN(n51) );
  AOI22_X1 U71 ( .A1(N115), .A2(n52), .B1(n51), .B2(n986), .ZN(n68) );
  AOI22_X1 U72 ( .A1(cta_id_mask_rev[12]), .A2(n59), .B1(cta_id_mask_rev[13]), 
        .B2(n58), .ZN(n53) );
  AOI221_X1 U73 ( .B1(cta_id_mask_rev[14]), .B2(n62), .C1(cta_id_mask_rev[15]), 
        .C2(n61), .A(n73), .ZN(n56) );
  AOI22_X1 U74 ( .A1(cta_id_mask_rev[8]), .A2(n59), .B1(cta_id_mask_rev[9]), 
        .B2(n58), .ZN(n54) );
  AOI221_X1 U75 ( .B1(cta_id_mask_rev[10]), .B2(n62), .C1(cta_id_mask_rev[11]), 
        .C2(n61), .A(n74), .ZN(n55) );
  OAI22_X1 U76 ( .A1(n987), .A2(n56), .B1(N114), .B2(n55), .ZN(n66) );
  AOI22_X1 U77 ( .A1(cta_id_mask_rev[4]), .A2(n59), .B1(cta_id_mask_rev[5]), 
        .B2(n58), .ZN(n57) );
  AOI221_X1 U78 ( .B1(cta_id_mask_rev[6]), .B2(n62), .C1(cta_id_mask_rev[7]), 
        .C2(n61), .A(n75), .ZN(n64) );
  AOI22_X1 U79 ( .A1(cta_id_mask_rev[0]), .A2(n59), .B1(cta_id_mask_rev[1]), 
        .B2(n58), .ZN(n60) );
  AOI221_X1 U80 ( .B1(cta_id_mask_rev[2]), .B2(n62), .C1(cta_id_mask_rev[3]), 
        .C2(n61), .A(n76), .ZN(n63) );
  OAI22_X1 U81 ( .A1(n987), .A2(n64), .B1(N114), .B2(n63), .ZN(n65) );
  AOI22_X1 U82 ( .A1(n66), .A2(N115), .B1(n65), .B2(n986), .ZN(n67) );
  OAI22_X1 U83 ( .A1(n68), .A2(n985), .B1(N116), .B2(n67), .ZN(N572) );
  INV_X1 U84 ( .A(n1), .ZN(n77) );
  INV_X1 U85 ( .A(n1), .ZN(n78) );
  INV_X1 U86 ( .A(n1), .ZN(n80) );
  INV_X1 U87 ( .A(n1), .ZN(n81) );
  CLKBUF_X1 U88 ( .A(n136), .Z(n109) );
  CLKBUF_X1 U89 ( .A(n136), .Z(n110) );
  CLKBUF_X1 U90 ( .A(n136), .Z(n111) );
  CLKBUF_X1 U91 ( .A(n136), .Z(n112) );
  CLKBUF_X1 U92 ( .A(n136), .Z(n113) );
  CLKBUF_X1 U93 ( .A(n136), .Z(n114) );
  CLKBUF_X1 U94 ( .A(n135), .Z(n115) );
  CLKBUF_X1 U95 ( .A(n135), .Z(n116) );
  CLKBUF_X1 U96 ( .A(n135), .Z(n117) );
  CLKBUF_X1 U97 ( .A(n135), .Z(n118) );
  CLKBUF_X1 U98 ( .A(n135), .Z(n119) );
  CLKBUF_X1 U99 ( .A(n135), .Z(n120) );
  CLKBUF_X1 U100 ( .A(n134), .Z(n121) );
  CLKBUF_X1 U101 ( .A(n134), .Z(n122) );
  CLKBUF_X1 U102 ( .A(n134), .Z(n123) );
  CLKBUF_X1 U103 ( .A(n134), .Z(n124) );
  CLKBUF_X1 U104 ( .A(n134), .Z(n125) );
  CLKBUF_X1 U105 ( .A(n134), .Z(n126) );
  CLKBUF_X1 U106 ( .A(n133), .Z(n127) );
  CLKBUF_X1 U107 ( .A(n133), .Z(n128) );
  CLKBUF_X1 U108 ( .A(n133), .Z(n129) );
  CLKBUF_X1 U109 ( .A(n133), .Z(n130) );
  CLKBUF_X1 U110 ( .A(n133), .Z(n131) );
  CLKBUF_X1 U111 ( .A(n133), .Z(n132) );
  XOR2_X1 U112 ( .A(\add_154/carry[5] ), .B(\warp_cntr[5] ), .Z(N707) );
  OAI221_X1 U113 ( .B1(n3), .B2(n145), .C1(n146), .C2(n147), .A(n148), .ZN(
        n651) );
  OAI22_X1 U114 ( .A1(n82), .A2(n807), .B1(n88), .B2(n150), .ZN(n999) );
  INV_X1 U115 ( .A(shmem_base_addr_in[4]), .ZN(n150) );
  OAI22_X1 U116 ( .A1(n79), .A2(n806), .B1(n83), .B2(n151), .ZN(n998) );
  INV_X1 U117 ( .A(shmem_base_addr_in[5]), .ZN(n151) );
  OAI22_X1 U118 ( .A1(n81), .A2(n805), .B1(n83), .B2(n152), .ZN(n997) );
  INV_X1 U119 ( .A(shmem_base_addr_in[6]), .ZN(n152) );
  OAI22_X1 U120 ( .A1(n80), .A2(n804), .B1(n83), .B2(n153), .ZN(n996) );
  INV_X1 U121 ( .A(shmem_base_addr_in[7]), .ZN(n153) );
  OAI22_X1 U122 ( .A1(n82), .A2(n803), .B1(n83), .B2(n154), .ZN(n995) );
  INV_X1 U123 ( .A(shmem_base_addr_in[8]), .ZN(n154) );
  OAI22_X1 U124 ( .A1(n82), .A2(n802), .B1(n83), .B2(n155), .ZN(n994) );
  INV_X1 U125 ( .A(shmem_base_addr_in[9]), .ZN(n155) );
  OAI22_X1 U126 ( .A1(n78), .A2(n801), .B1(n83), .B2(n156), .ZN(n993) );
  INV_X1 U127 ( .A(shmem_base_addr_in[10]), .ZN(n156) );
  OAI22_X1 U128 ( .A1(n77), .A2(n800), .B1(n83), .B2(n157), .ZN(n992) );
  INV_X1 U129 ( .A(shmem_base_addr_in[11]), .ZN(n157) );
  OAI22_X1 U130 ( .A1(n82), .A2(n799), .B1(n84), .B2(n158), .ZN(n991) );
  INV_X1 U131 ( .A(shmem_base_addr_in[12]), .ZN(n158) );
  OAI22_X1 U132 ( .A1(n79), .A2(n798), .B1(n83), .B2(n159), .ZN(n990) );
  INV_X1 U133 ( .A(shmem_base_addr_in[13]), .ZN(n159) );
  OAI22_X1 U134 ( .A1(n160), .A2(n917), .B1(n161), .B2(n162), .ZN(n984) );
  OAI21_X1 U135 ( .B1(n9), .B2(n96), .A(n164), .ZN(n983) );
  NAND2_X1 U136 ( .A1(N707), .A2(n165), .ZN(n164) );
  NOR2_X1 U137 ( .A1(reset), .A2(host_reset), .ZN(n982) );
  OAI21_X1 U138 ( .B1(n166), .B2(n167), .A(n10), .ZN(n981) );
  OAI21_X1 U139 ( .B1(n166), .B2(n168), .A(n11), .ZN(n980) );
  OAI21_X1 U140 ( .B1(n166), .B2(n169), .A(n12), .ZN(n979) );
  OAI21_X1 U141 ( .B1(n166), .B2(n170), .A(n13), .ZN(n978) );
  OAI21_X1 U142 ( .B1(n166), .B2(n171), .A(n14), .ZN(n977) );
  OAI21_X1 U143 ( .B1(n166), .B2(n172), .A(n15), .ZN(n976) );
  OAI21_X1 U144 ( .B1(n166), .B2(n173), .A(n16), .ZN(n975) );
  OAI21_X1 U145 ( .B1(n166), .B2(n174), .A(n17), .ZN(n974) );
  NAND3_X1 U146 ( .A1(warp_id_in[3]), .A2(n175), .A3(warp_id_in[4]), .ZN(n166)
         );
  OAI21_X1 U147 ( .B1(n167), .B2(n176), .A(n18), .ZN(n973) );
  OAI21_X1 U148 ( .B1(n168), .B2(n176), .A(n19), .ZN(n972) );
  OAI21_X1 U149 ( .B1(n169), .B2(n176), .A(n20), .ZN(n971) );
  OAI21_X1 U150 ( .B1(n170), .B2(n176), .A(n21), .ZN(n970) );
  OAI21_X1 U151 ( .B1(n171), .B2(n176), .A(n22), .ZN(n969) );
  OAI21_X1 U152 ( .B1(n172), .B2(n176), .A(n23), .ZN(n968) );
  OAI21_X1 U153 ( .B1(n173), .B2(n176), .A(n24), .ZN(n967) );
  OAI21_X1 U154 ( .B1(n174), .B2(n176), .A(n25), .ZN(n966) );
  NAND3_X1 U155 ( .A1(n175), .A2(n177), .A3(warp_id_in[4]), .ZN(n176) );
  OAI21_X1 U156 ( .B1(n167), .B2(n178), .A(n26), .ZN(n965) );
  OAI21_X1 U157 ( .B1(n168), .B2(n178), .A(n27), .ZN(n964) );
  OAI21_X1 U158 ( .B1(n169), .B2(n178), .A(n28), .ZN(n963) );
  OAI21_X1 U159 ( .B1(n170), .B2(n178), .A(n29), .ZN(n962) );
  OAI21_X1 U160 ( .B1(n171), .B2(n178), .A(n30), .ZN(n961) );
  OAI21_X1 U161 ( .B1(n172), .B2(n178), .A(n31), .ZN(n960) );
  OAI21_X1 U162 ( .B1(n173), .B2(n178), .A(n32), .ZN(n959) );
  OAI21_X1 U163 ( .B1(n174), .B2(n178), .A(n33), .ZN(n958) );
  NAND3_X1 U164 ( .A1(n175), .A2(n179), .A3(warp_id_in[3]), .ZN(n178) );
  OAI21_X1 U165 ( .B1(n167), .B2(n180), .A(n34), .ZN(n957) );
  OAI21_X1 U166 ( .B1(n168), .B2(n180), .A(n35), .ZN(n956) );
  OAI21_X1 U167 ( .B1(n169), .B2(n180), .A(n36), .ZN(n955) );
  OAI21_X1 U168 ( .B1(n170), .B2(n180), .A(n37), .ZN(n954) );
  OAI21_X1 U169 ( .B1(n171), .B2(n180), .A(n38), .ZN(n953) );
  OAI21_X1 U170 ( .B1(n172), .B2(n180), .A(n39), .ZN(n952) );
  OAI21_X1 U171 ( .B1(n173), .B2(n180), .A(n40), .ZN(n951) );
  OAI21_X1 U172 ( .B1(n174), .B2(n180), .A(n41), .ZN(n950) );
  NAND3_X1 U173 ( .A1(n177), .A2(n179), .A3(n175), .ZN(n180) );
  AND4_X1 U174 ( .A1(warp_state_in[0]), .A2(n181), .A3(warp_state_in[1]), .A4(
        n182), .ZN(n175) );
  MUX2_X1 U175 ( .A(warp_checker_state_machine[2]), .B(n183), .S(n145), .Z(
        n1267) );
  OAI221_X1 U176 ( .B1(N567), .B2(n146), .C1(n184), .C2(n185), .A(n186), .ZN(
        n183) );
  OAI221_X1 U177 ( .B1(n7), .B2(n145), .C1(n146), .C2(n147), .A(n187), .ZN(
        n1266) );
  INV_X1 U178 ( .A(N567), .ZN(n147) );
  NAND4_X1 U179 ( .A1(n102), .A2(n187), .A3(n146), .A4(n188), .ZN(n145) );
  AOI21_X1 U180 ( .B1(\warp_cntr[5] ), .B2(n189), .A(n190), .ZN(n188) );
  NAND3_X1 U181 ( .A1(n3), .A2(n8), .A3(warp_checker_state_machine[1]), .ZN(
        n146) );
  OAI21_X1 U182 ( .B1(n988), .B2(n96), .A(n191), .ZN(n1265) );
  NAND2_X1 U183 ( .A1(N703), .A2(n165), .ZN(n191) );
  OAI21_X1 U184 ( .B1(n989), .B2(n96), .A(n192), .ZN(n1264) );
  NAND2_X1 U185 ( .A1(n989), .A2(n165), .ZN(n192) );
  OAI21_X1 U186 ( .B1(n987), .B2(n96), .A(n193), .ZN(n1263) );
  NAND2_X1 U187 ( .A1(N704), .A2(n165), .ZN(n193) );
  OAI21_X1 U188 ( .B1(n986), .B2(n96), .A(n194), .ZN(n1262) );
  NAND2_X1 U189 ( .A1(N705), .A2(n165), .ZN(n194) );
  OAI21_X1 U190 ( .B1(n985), .B2(n96), .A(n195), .ZN(n1261) );
  NAND2_X1 U191 ( .A1(N706), .A2(n165), .ZN(n195) );
  MUX2_X1 U192 ( .A(warp_id_in[0]), .B(warp_id_addr[0]), .S(n101), .Z(n1260)
         );
  MUX2_X1 U193 ( .A(warp_id_in[4]), .B(warp_id_addr[4]), .S(n101), .Z(n1259)
         );
  MUX2_X1 U194 ( .A(warp_id_in[3]), .B(warp_id_addr[3]), .S(n101), .Z(n1258)
         );
  MUX2_X1 U195 ( .A(warp_id_in[2]), .B(warp_id_addr[2]), .S(n101), .Z(n1257)
         );
  MUX2_X1 U196 ( .A(warp_id_in[1]), .B(warp_id_addr[1]), .S(n101), .Z(n1256)
         );
  NAND2_X1 U197 ( .A1(n185), .A2(n196), .ZN(n1255) );
  NAND3_X1 U198 ( .A1(n197), .A2(n102), .A3(pipeline_stall_out), .ZN(n196) );
  INV_X1 U199 ( .A(n181), .ZN(n185) );
  MUX2_X1 U200 ( .A(n96), .B(fence_regs_fence_en_ld[0]), .S(n198), .Z(n1254)
         );
  AOI21_X1 U201 ( .B1(n199), .B2(n200), .A(n201), .ZN(n198) );
  MUX2_X1 U202 ( .A(n96), .B(fence_regs_fence_en_ld[1]), .S(n202), .Z(n1253)
         );
  AOI21_X1 U203 ( .B1(n203), .B2(n200), .A(n204), .ZN(n202) );
  MUX2_X1 U204 ( .A(n96), .B(fence_regs_fence_en_ld[2]), .S(n205), .Z(n1252)
         );
  AOI21_X1 U205 ( .B1(n206), .B2(n200), .A(n207), .ZN(n205) );
  MUX2_X1 U206 ( .A(n96), .B(fence_regs_fence_en_ld[3]), .S(n208), .Z(n1251)
         );
  AOI21_X1 U207 ( .B1(n209), .B2(n200), .A(n210), .ZN(n208) );
  MUX2_X1 U208 ( .A(n96), .B(fence_regs_fence_en_ld[4]), .S(n211), .Z(n1250)
         );
  AOI21_X1 U209 ( .B1(n212), .B2(n200), .A(n213), .ZN(n211) );
  MUX2_X1 U210 ( .A(n96), .B(fence_regs_fence_en_ld[5]), .S(n214), .Z(n1249)
         );
  AOI21_X1 U211 ( .B1(n215), .B2(n200), .A(n216), .ZN(n214) );
  MUX2_X1 U212 ( .A(n96), .B(fence_regs_fence_en_ld[6]), .S(n217), .Z(n1248)
         );
  AOI21_X1 U213 ( .B1(n218), .B2(n200), .A(n219), .ZN(n217) );
  MUX2_X1 U214 ( .A(n96), .B(fence_regs_fence_en_ld[7]), .S(n220), .Z(n1247)
         );
  AOI21_X1 U215 ( .B1(n221), .B2(n200), .A(n222), .ZN(n220) );
  MUX2_X1 U216 ( .A(n97), .B(fence_regs_fence_en_ld[8]), .S(n223), .Z(n1246)
         );
  AOI21_X1 U217 ( .B1(n224), .B2(n199), .A(n225), .ZN(n223) );
  MUX2_X1 U218 ( .A(n97), .B(fence_regs_fence_en_ld[9]), .S(n226), .Z(n1245)
         );
  AOI21_X1 U219 ( .B1(n224), .B2(n203), .A(n227), .ZN(n226) );
  MUX2_X1 U220 ( .A(n97), .B(fence_regs_fence_en_ld[10]), .S(n228), .Z(n1244)
         );
  AOI21_X1 U221 ( .B1(n224), .B2(n206), .A(n229), .ZN(n228) );
  MUX2_X1 U222 ( .A(n97), .B(fence_regs_fence_en_ld[11]), .S(n230), .Z(n1243)
         );
  AOI21_X1 U223 ( .B1(n224), .B2(n209), .A(n231), .ZN(n230) );
  MUX2_X1 U224 ( .A(n97), .B(fence_regs_fence_en_ld[12]), .S(n232), .Z(n1242)
         );
  AOI21_X1 U225 ( .B1(n224), .B2(n212), .A(n233), .ZN(n232) );
  MUX2_X1 U226 ( .A(n97), .B(fence_regs_fence_en_ld[13]), .S(n234), .Z(n1241)
         );
  AOI21_X1 U227 ( .B1(n224), .B2(n215), .A(n235), .ZN(n234) );
  MUX2_X1 U228 ( .A(n97), .B(fence_regs_fence_en_ld[14]), .S(n236), .Z(n1240)
         );
  AOI21_X1 U229 ( .B1(n224), .B2(n218), .A(n237), .ZN(n236) );
  MUX2_X1 U230 ( .A(n97), .B(fence_regs_fence_en_ld[15]), .S(n238), .Z(n1239)
         );
  AOI21_X1 U231 ( .B1(n224), .B2(n221), .A(n239), .ZN(n238) );
  MUX2_X1 U232 ( .A(n97), .B(fence_regs_fence_en_ld[16]), .S(n240), .Z(n1238)
         );
  AOI21_X1 U233 ( .B1(n241), .B2(n199), .A(n242), .ZN(n240) );
  MUX2_X1 U234 ( .A(n97), .B(fence_regs_fence_en_ld[17]), .S(n243), .Z(n1237)
         );
  AOI21_X1 U235 ( .B1(n241), .B2(n203), .A(n244), .ZN(n243) );
  MUX2_X1 U236 ( .A(n97), .B(fence_regs_fence_en_ld[18]), .S(n245), .Z(n1236)
         );
  AOI21_X1 U237 ( .B1(n241), .B2(n206), .A(n246), .ZN(n245) );
  MUX2_X1 U238 ( .A(n97), .B(fence_regs_fence_en_ld[19]), .S(n247), .Z(n1235)
         );
  AOI21_X1 U239 ( .B1(n241), .B2(n209), .A(n248), .ZN(n247) );
  MUX2_X1 U240 ( .A(n97), .B(fence_regs_fence_en_ld[20]), .S(n249), .Z(n1234)
         );
  AOI21_X1 U241 ( .B1(n241), .B2(n212), .A(n250), .ZN(n249) );
  MUX2_X1 U242 ( .A(n97), .B(fence_regs_fence_en_ld[21]), .S(n251), .Z(n1233)
         );
  AOI21_X1 U243 ( .B1(n241), .B2(n215), .A(n252), .ZN(n251) );
  MUX2_X1 U244 ( .A(n97), .B(fence_regs_fence_en_ld[22]), .S(n253), .Z(n1232)
         );
  AOI21_X1 U245 ( .B1(n241), .B2(n218), .A(n254), .ZN(n253) );
  MUX2_X1 U246 ( .A(n97), .B(fence_regs_fence_en_ld[23]), .S(n255), .Z(n1231)
         );
  AOI21_X1 U247 ( .B1(n241), .B2(n221), .A(n256), .ZN(n255) );
  AND3_X1 U248 ( .A1(warp_id_addr[4]), .A2(n6), .A3(n257), .ZN(n241) );
  MUX2_X1 U249 ( .A(n98), .B(fence_regs_fence_en_ld[24]), .S(n258), .Z(n1230)
         );
  AOI21_X1 U250 ( .B1(n259), .B2(n199), .A(n260), .ZN(n258) );
  NOR3_X1 U251 ( .A1(warp_id_addr[1]), .A2(warp_id_addr[2]), .A3(
        warp_id_addr[0]), .ZN(n199) );
  MUX2_X1 U252 ( .A(n98), .B(fence_regs_fence_en_ld[25]), .S(n261), .Z(n1229)
         );
  AOI21_X1 U253 ( .B1(n259), .B2(n203), .A(n262), .ZN(n261) );
  NOR3_X1 U254 ( .A1(warp_id_addr[1]), .A2(warp_id_addr[2]), .A3(n4), .ZN(n203) );
  MUX2_X1 U255 ( .A(n98), .B(fence_regs_fence_en_ld[26]), .S(n263), .Z(n1228)
         );
  AOI21_X1 U256 ( .B1(n259), .B2(n206), .A(n264), .ZN(n263) );
  NOR3_X1 U257 ( .A1(warp_id_addr[0]), .A2(warp_id_addr[2]), .A3(n5), .ZN(n206) );
  MUX2_X1 U258 ( .A(n98), .B(fence_regs_fence_en_ld[27]), .S(n265), .Z(n1227)
         );
  AOI21_X1 U259 ( .B1(n259), .B2(n209), .A(n266), .ZN(n265) );
  NOR3_X1 U260 ( .A1(n4), .A2(warp_id_addr[2]), .A3(n5), .ZN(n209) );
  MUX2_X1 U261 ( .A(n98), .B(fence_regs_fence_en_ld[28]), .S(n267), .Z(n1226)
         );
  AOI21_X1 U262 ( .B1(n259), .B2(n212), .A(n268), .ZN(n267) );
  AND3_X1 U263 ( .A1(n4), .A2(n5), .A3(warp_id_addr[2]), .ZN(n212) );
  MUX2_X1 U264 ( .A(n98), .B(fence_regs_fence_en_ld[29]), .S(n269), .Z(n1225)
         );
  AOI21_X1 U265 ( .B1(n259), .B2(n215), .A(n270), .ZN(n269) );
  AND3_X1 U266 ( .A1(warp_id_addr[0]), .A2(n5), .A3(warp_id_addr[2]), .ZN(n215) );
  MUX2_X1 U267 ( .A(n98), .B(fence_regs_fence_en_ld[30]), .S(n271), .Z(n1224)
         );
  AOI21_X1 U268 ( .B1(n259), .B2(n218), .A(n272), .ZN(n271) );
  AND3_X1 U269 ( .A1(warp_id_addr[2]), .A2(n4), .A3(warp_id_addr[1]), .ZN(n218) );
  MUX2_X1 U270 ( .A(n98), .B(fence_regs_fence_en_ld[31]), .S(n273), .Z(n1223)
         );
  AOI21_X1 U271 ( .B1(n259), .B2(n221), .A(n274), .ZN(n273) );
  AND3_X1 U272 ( .A1(warp_id_addr[2]), .A2(warp_id_addr[0]), .A3(
        warp_id_addr[1]), .ZN(n221) );
  AND3_X1 U273 ( .A1(warp_id_addr[3]), .A2(warp_id_addr[4]), .A3(n257), .ZN(
        n259) );
  NAND2_X1 U274 ( .A1(n186), .A2(n102), .ZN(n163) );
  INV_X1 U275 ( .A(n189), .ZN(n186) );
  OAI22_X1 U276 ( .A1(n78), .A2(n781), .B1(n84), .B2(n275), .ZN(n1222) );
  OAI22_X1 U277 ( .A1(n77), .A2(n782), .B1(n83), .B2(n144), .ZN(n1221) );
  OAI22_X1 U278 ( .A1(n77), .A2(n783), .B1(n84), .B2(n142), .ZN(n1220) );
  OAI22_X1 U279 ( .A1(n77), .A2(n784), .B1(n84), .B2(n140), .ZN(n1219) );
  OAI22_X1 U280 ( .A1(n77), .A2(n785), .B1(n84), .B2(n138), .ZN(n1218) );
  OAI22_X1 U281 ( .A1(n77), .A2(n786), .B1(n84), .B2(n276), .ZN(n1217) );
  OAI21_X1 U282 ( .B1(n82), .B2(n787), .A(n83), .ZN(n1216) );
  OAI22_X1 U283 ( .A1(n77), .A2(n788), .B1(n84), .B2(n179), .ZN(n1215) );
  OAI22_X1 U284 ( .A1(n77), .A2(n789), .B1(n84), .B2(n177), .ZN(n1214) );
  OAI22_X1 U285 ( .A1(n77), .A2(n790), .B1(n84), .B2(n277), .ZN(n1213) );
  OAI222_X1 U286 ( .A1(n989), .A2(n278), .B1(n162), .B2(n275), .C1(n160), .C2(
        n791), .ZN(n1212) );
  OAI21_X1 U287 ( .B1(n160), .B2(n1173), .A(n279), .ZN(n1211) );
  NAND3_X1 U288 ( .A1(n280), .A2(warp_state_in[1]), .A3(warp_state_in[0]), 
        .ZN(n279) );
  INV_X1 U289 ( .A(n162), .ZN(n280) );
  OAI222_X1 U290 ( .A1(n985), .A2(n278), .B1(n162), .B2(n179), .C1(n160), .C2(
        n792), .ZN(n1210) );
  OAI222_X1 U291 ( .A1(n986), .A2(n278), .B1(n162), .B2(n177), .C1(n160), .C2(
        n793), .ZN(n1209) );
  OAI222_X1 U292 ( .A1(n987), .A2(n278), .B1(n162), .B2(n277), .C1(n160), .C2(
        n794), .ZN(n1208) );
  OAI222_X1 U293 ( .A1(n988), .A2(n278), .B1(n162), .B2(n276), .C1(n160), .C2(
        n795), .ZN(n1207) );
  NAND2_X1 U294 ( .A1(n181), .A2(n160), .ZN(n162) );
  NAND2_X1 U295 ( .A1(n189), .A2(n160), .ZN(n278) );
  OAI211_X1 U296 ( .C1(n796), .C2(n282), .A(n281), .B(n83), .ZN(n1206) );
  NAND2_X1 U297 ( .A1(n1), .A2(n283), .ZN(n282) );
  MUX2_X1 U298 ( .A(fence_regs_fence_en_out[0]), .B(n100), .S(n201), .Z(n1205)
         );
  OAI22_X1 U299 ( .A1(n174), .A2(n284), .B1(n285), .B2(n286), .ZN(n201) );
  MUX2_X1 U300 ( .A(fence_regs_fence_en_out[31]), .B(n100), .S(n274), .Z(n1204) );
  OAI22_X1 U301 ( .A1(n167), .A2(n287), .B1(n288), .B2(n289), .ZN(n274) );
  MUX2_X1 U302 ( .A(fence_regs_fence_en_out[30]), .B(n100), .S(n272), .Z(n1203) );
  OAI22_X1 U303 ( .A1(n168), .A2(n287), .B1(n290), .B2(n289), .ZN(n272) );
  MUX2_X1 U304 ( .A(fence_regs_fence_en_out[29]), .B(n100), .S(n270), .Z(n1202) );
  OAI22_X1 U305 ( .A1(n169), .A2(n287), .B1(n291), .B2(n289), .ZN(n270) );
  MUX2_X1 U306 ( .A(fence_regs_fence_en_out[28]), .B(n100), .S(n268), .Z(n1201) );
  OAI22_X1 U307 ( .A1(n170), .A2(n287), .B1(n292), .B2(n289), .ZN(n268) );
  MUX2_X1 U308 ( .A(fence_regs_fence_en_out[27]), .B(n100), .S(n266), .Z(n1200) );
  OAI22_X1 U309 ( .A1(n171), .A2(n287), .B1(n293), .B2(n289), .ZN(n266) );
  MUX2_X1 U310 ( .A(fence_regs_fence_en_out[26]), .B(n100), .S(n264), .Z(n1199) );
  OAI22_X1 U311 ( .A1(n172), .A2(n287), .B1(n294), .B2(n289), .ZN(n264) );
  MUX2_X1 U312 ( .A(fence_regs_fence_en_out[25]), .B(n100), .S(n262), .Z(n1198) );
  OAI22_X1 U313 ( .A1(n173), .A2(n287), .B1(n295), .B2(n289), .ZN(n262) );
  MUX2_X1 U314 ( .A(fence_regs_fence_en_out[24]), .B(n100), .S(n260), .Z(n1197) );
  OAI22_X1 U315 ( .A1(n174), .A2(n287), .B1(n285), .B2(n289), .ZN(n260) );
  NAND3_X1 U316 ( .A1(N116), .A2(N115), .A3(n296), .ZN(n289) );
  NAND3_X1 U317 ( .A1(warp_id_in[4]), .A2(warp_id_in[3]), .A3(n297), .ZN(n287)
         );
  MUX2_X1 U318 ( .A(fence_regs_fence_en_out[23]), .B(n100), .S(n256), .Z(n1196) );
  OAI22_X1 U319 ( .A1(n167), .A2(n298), .B1(n288), .B2(n299), .ZN(n256) );
  MUX2_X1 U320 ( .A(fence_regs_fence_en_out[22]), .B(n100), .S(n254), .Z(n1195) );
  OAI22_X1 U321 ( .A1(n168), .A2(n298), .B1(n290), .B2(n299), .ZN(n254) );
  MUX2_X1 U322 ( .A(fence_regs_fence_en_out[21]), .B(n100), .S(n252), .Z(n1194) );
  OAI22_X1 U323 ( .A1(n169), .A2(n298), .B1(n291), .B2(n299), .ZN(n252) );
  MUX2_X1 U324 ( .A(fence_regs_fence_en_out[20]), .B(n100), .S(n250), .Z(n1193) );
  OAI22_X1 U325 ( .A1(n170), .A2(n298), .B1(n292), .B2(n299), .ZN(n250) );
  MUX2_X1 U326 ( .A(fence_regs_fence_en_out[19]), .B(n100), .S(n248), .Z(n1192) );
  OAI22_X1 U327 ( .A1(n171), .A2(n298), .B1(n293), .B2(n299), .ZN(n248) );
  MUX2_X1 U328 ( .A(fence_regs_fence_en_out[18]), .B(n100), .S(n246), .Z(n1191) );
  OAI22_X1 U329 ( .A1(n172), .A2(n298), .B1(n294), .B2(n299), .ZN(n246) );
  MUX2_X1 U330 ( .A(fence_regs_fence_en_out[17]), .B(n100), .S(n244), .Z(n1190) );
  OAI22_X1 U331 ( .A1(n173), .A2(n298), .B1(n295), .B2(n299), .ZN(n244) );
  MUX2_X1 U332 ( .A(fence_regs_fence_en_out[16]), .B(n100), .S(n242), .Z(n1189) );
  OAI22_X1 U333 ( .A1(n174), .A2(n298), .B1(n285), .B2(n299), .ZN(n242) );
  NAND3_X1 U334 ( .A1(n296), .A2(N116), .A3(n986), .ZN(n299) );
  NAND3_X1 U335 ( .A1(warp_id_in[4]), .A2(n177), .A3(n297), .ZN(n298) );
  MUX2_X1 U336 ( .A(fence_regs_fence_en_out[15]), .B(n100), .S(n239), .Z(n1188) );
  OAI22_X1 U337 ( .A1(n167), .A2(n300), .B1(n288), .B2(n301), .ZN(n239) );
  MUX2_X1 U338 ( .A(fence_regs_fence_en_out[14]), .B(n99), .S(n237), .Z(n1187)
         );
  OAI22_X1 U339 ( .A1(n168), .A2(n300), .B1(n290), .B2(n301), .ZN(n237) );
  MUX2_X1 U340 ( .A(fence_regs_fence_en_out[13]), .B(n99), .S(n235), .Z(n1186)
         );
  OAI22_X1 U341 ( .A1(n169), .A2(n300), .B1(n291), .B2(n301), .ZN(n235) );
  MUX2_X1 U342 ( .A(fence_regs_fence_en_out[12]), .B(n99), .S(n233), .Z(n1185)
         );
  OAI22_X1 U343 ( .A1(n170), .A2(n300), .B1(n292), .B2(n301), .ZN(n233) );
  MUX2_X1 U344 ( .A(fence_regs_fence_en_out[11]), .B(n99), .S(n231), .Z(n1184)
         );
  OAI22_X1 U345 ( .A1(n171), .A2(n300), .B1(n293), .B2(n301), .ZN(n231) );
  MUX2_X1 U346 ( .A(fence_regs_fence_en_out[10]), .B(n99), .S(n229), .Z(n1183)
         );
  OAI22_X1 U347 ( .A1(n172), .A2(n300), .B1(n294), .B2(n301), .ZN(n229) );
  MUX2_X1 U348 ( .A(fence_regs_fence_en_out[9]), .B(n99), .S(n227), .Z(n1182)
         );
  OAI22_X1 U349 ( .A1(n173), .A2(n300), .B1(n295), .B2(n301), .ZN(n227) );
  MUX2_X1 U350 ( .A(fence_regs_fence_en_out[8]), .B(n99), .S(n225), .Z(n1181)
         );
  OAI22_X1 U351 ( .A1(n174), .A2(n300), .B1(n285), .B2(n301), .ZN(n225) );
  NAND3_X1 U352 ( .A1(n296), .A2(N115), .A3(n985), .ZN(n301) );
  NAND3_X1 U353 ( .A1(n988), .A2(n987), .A3(n989), .ZN(n285) );
  NAND3_X1 U354 ( .A1(warp_id_in[3]), .A2(n179), .A3(n297), .ZN(n300) );
  NAND3_X1 U355 ( .A1(n276), .A2(n277), .A3(n275), .ZN(n174) );
  MUX2_X1 U356 ( .A(fence_regs_fence_en_out[7]), .B(n99), .S(n222), .Z(n1180)
         );
  OAI22_X1 U357 ( .A1(n167), .A2(n284), .B1(n286), .B2(n288), .ZN(n222) );
  NAND3_X1 U358 ( .A1(N113), .A2(N112), .A3(N114), .ZN(n288) );
  NAND3_X1 U359 ( .A1(warp_id_in[1]), .A2(warp_id_in[0]), .A3(warp_id_in[2]), 
        .ZN(n167) );
  MUX2_X1 U360 ( .A(fence_regs_fence_en_out[6]), .B(n99), .S(n219), .Z(n1179)
         );
  OAI22_X1 U361 ( .A1(n168), .A2(n284), .B1(n286), .B2(n290), .ZN(n219) );
  NAND3_X1 U362 ( .A1(N114), .A2(N113), .A3(n989), .ZN(n290) );
  NAND3_X1 U363 ( .A1(warp_id_in[1]), .A2(n275), .A3(warp_id_in[2]), .ZN(n168)
         );
  MUX2_X1 U364 ( .A(fence_regs_fence_en_out[5]), .B(n99), .S(n216), .Z(n1178)
         );
  OAI22_X1 U365 ( .A1(n169), .A2(n284), .B1(n286), .B2(n291), .ZN(n216) );
  NAND3_X1 U366 ( .A1(N114), .A2(N112), .A3(n988), .ZN(n291) );
  NAND3_X1 U367 ( .A1(warp_id_in[0]), .A2(n276), .A3(warp_id_in[2]), .ZN(n169)
         );
  MUX2_X1 U368 ( .A(fence_regs_fence_en_out[4]), .B(n99), .S(n213), .Z(n1177)
         );
  OAI22_X1 U369 ( .A1(n170), .A2(n284), .B1(n286), .B2(n292), .ZN(n213) );
  NAND3_X1 U370 ( .A1(n988), .A2(N114), .A3(n989), .ZN(n292) );
  NAND3_X1 U371 ( .A1(n275), .A2(n276), .A3(warp_id_in[2]), .ZN(n170) );
  MUX2_X1 U372 ( .A(fence_regs_fence_en_out[3]), .B(n99), .S(n210), .Z(n1176)
         );
  OAI22_X1 U373 ( .A1(n171), .A2(n284), .B1(n286), .B2(n293), .ZN(n210) );
  NAND3_X1 U374 ( .A1(N113), .A2(N112), .A3(n987), .ZN(n293) );
  NAND3_X1 U375 ( .A1(warp_id_in[0]), .A2(n277), .A3(warp_id_in[1]), .ZN(n171)
         );
  MUX2_X1 U376 ( .A(fence_regs_fence_en_out[2]), .B(n99), .S(n207), .Z(n1175)
         );
  OAI22_X1 U377 ( .A1(n172), .A2(n284), .B1(n286), .B2(n294), .ZN(n207) );
  NAND3_X1 U378 ( .A1(n987), .A2(N113), .A3(n989), .ZN(n294) );
  NAND3_X1 U379 ( .A1(n275), .A2(n277), .A3(warp_id_in[1]), .ZN(n172) );
  INV_X1 U380 ( .A(warp_id_in[0]), .ZN(n275) );
  MUX2_X1 U381 ( .A(fence_regs_fence_en_out[1]), .B(n99), .S(n204), .Z(n1174)
         );
  OAI22_X1 U382 ( .A1(n173), .A2(n284), .B1(n286), .B2(n295), .ZN(n204) );
  NAND3_X1 U383 ( .A1(n987), .A2(N112), .A3(n988), .ZN(n295) );
  NAND3_X1 U384 ( .A1(n985), .A2(n296), .A3(n986), .ZN(n286) );
  INV_X1 U385 ( .A(n281), .ZN(n296) );
  NAND2_X1 U386 ( .A1(N572), .A2(n165), .ZN(n281) );
  INV_X1 U387 ( .A(n283), .ZN(n165) );
  NAND2_X1 U388 ( .A1(n9), .A2(n189), .ZN(n283) );
  NOR3_X1 U389 ( .A1(n3), .A2(warp_checker_state_machine[2]), .A3(n7), .ZN(
        n189) );
  NAND3_X1 U390 ( .A1(n177), .A2(n179), .A3(n297), .ZN(n284) );
  INV_X1 U391 ( .A(n148), .ZN(n297) );
  NAND2_X1 U392 ( .A1(n181), .A2(n184), .ZN(n148) );
  NOR3_X1 U393 ( .A1(n302), .A2(warp_state_in[0]), .A3(n161), .ZN(n184) );
  INV_X1 U394 ( .A(warp_state_in[1]), .ZN(n161) );
  INV_X1 U395 ( .A(warp_id_in[4]), .ZN(n179) );
  INV_X1 U396 ( .A(warp_id_in[3]), .ZN(n177) );
  NAND3_X1 U397 ( .A1(n276), .A2(n277), .A3(warp_id_in[0]), .ZN(n173) );
  INV_X1 U398 ( .A(warp_id_in[2]), .ZN(n277) );
  INV_X1 U399 ( .A(warp_id_in[1]), .ZN(n276) );
  MUX2_X1 U400 ( .A(warps_done_mask[0]), .B(warps_done_mask_out[0]), .S(n106), 
        .Z(n1140) );
  MUX2_X1 U401 ( .A(warps_done_mask[1]), .B(warps_done_mask_out[1]), .S(n106), 
        .Z(n1139) );
  MUX2_X1 U402 ( .A(warps_done_mask[2]), .B(warps_done_mask_out[2]), .S(n106), 
        .Z(n1138) );
  MUX2_X1 U403 ( .A(warps_done_mask[3]), .B(warps_done_mask_out[3]), .S(n106), 
        .Z(n1137) );
  MUX2_X1 U404 ( .A(warps_done_mask[4]), .B(warps_done_mask_out[4]), .S(n106), 
        .Z(n1136) );
  MUX2_X1 U405 ( .A(warps_done_mask[5]), .B(warps_done_mask_out[5]), .S(n106), 
        .Z(n1135) );
  MUX2_X1 U406 ( .A(warps_done_mask[6]), .B(warps_done_mask_out[6]), .S(n106), 
        .Z(n1134) );
  MUX2_X1 U407 ( .A(warps_done_mask[7]), .B(warps_done_mask_out[7]), .S(n106), 
        .Z(n1133) );
  MUX2_X1 U408 ( .A(warps_done_mask[8]), .B(warps_done_mask_out[8]), .S(n105), 
        .Z(n1132) );
  MUX2_X1 U409 ( .A(warps_done_mask[9]), .B(warps_done_mask_out[9]), .S(n105), 
        .Z(n1131) );
  MUX2_X1 U410 ( .A(warps_done_mask[10]), .B(warps_done_mask_out[10]), .S(n105), .Z(n1130) );
  MUX2_X1 U411 ( .A(warps_done_mask[11]), .B(warps_done_mask_out[11]), .S(n105), .Z(n1129) );
  MUX2_X1 U412 ( .A(warps_done_mask[12]), .B(warps_done_mask_out[12]), .S(n105), .Z(n1128) );
  MUX2_X1 U413 ( .A(warps_done_mask[13]), .B(warps_done_mask_out[13]), .S(n105), .Z(n1127) );
  MUX2_X1 U414 ( .A(warps_done_mask[14]), .B(warps_done_mask_out[14]), .S(n105), .Z(n1126) );
  MUX2_X1 U415 ( .A(warps_done_mask[15]), .B(warps_done_mask_out[15]), .S(n105), .Z(n1125) );
  MUX2_X1 U416 ( .A(warps_done_mask[16]), .B(warps_done_mask_out[16]), .S(n105), .Z(n1124) );
  MUX2_X1 U417 ( .A(warps_done_mask[17]), .B(warps_done_mask_out[17]), .S(n105), .Z(n1123) );
  MUX2_X1 U418 ( .A(warps_done_mask[18]), .B(warps_done_mask_out[18]), .S(n105), .Z(n1122) );
  MUX2_X1 U419 ( .A(warps_done_mask[19]), .B(warps_done_mask_out[19]), .S(n105), .Z(n1121) );
  MUX2_X1 U420 ( .A(warps_done_mask[20]), .B(warps_done_mask_out[20]), .S(n104), .Z(n1120) );
  MUX2_X1 U421 ( .A(warps_done_mask[21]), .B(warps_done_mask_out[21]), .S(n104), .Z(n1119) );
  MUX2_X1 U422 ( .A(warps_done_mask[22]), .B(warps_done_mask_out[22]), .S(n104), .Z(n1118) );
  MUX2_X1 U423 ( .A(warps_done_mask[23]), .B(warps_done_mask_out[23]), .S(n104), .Z(n1117) );
  MUX2_X1 U424 ( .A(warps_done_mask[24]), .B(warps_done_mask_out[24]), .S(n104), .Z(n1116) );
  MUX2_X1 U425 ( .A(warps_done_mask[25]), .B(warps_done_mask_out[25]), .S(n104), .Z(n1115) );
  MUX2_X1 U426 ( .A(warps_done_mask[26]), .B(warps_done_mask_out[26]), .S(n104), .Z(n1114) );
  MUX2_X1 U427 ( .A(warps_done_mask[27]), .B(warps_done_mask_out[27]), .S(n104), .Z(n1113) );
  MUX2_X1 U428 ( .A(warps_done_mask[28]), .B(warps_done_mask_out[28]), .S(n104), .Z(n1112) );
  MUX2_X1 U429 ( .A(warps_done_mask[29]), .B(warps_done_mask_out[29]), .S(n104), .Z(n1111) );
  MUX2_X1 U430 ( .A(warps_done_mask[30]), .B(warps_done_mask_out[30]), .S(n104), .Z(n1110) );
  MUX2_X1 U431 ( .A(warps_done_mask[31]), .B(warps_done_mask_out[31]), .S(n104), .Z(n1109) );
  AOI21_X1 U432 ( .B1(n304), .B2(n99), .A(n190), .ZN(n303) );
  OAI22_X1 U433 ( .A1(n77), .A2(n916), .B1(n84), .B2(n305), .ZN(n1108) );
  INV_X1 U434 ( .A(current_mask_in[0]), .ZN(n305) );
  OAI22_X1 U435 ( .A1(n77), .A2(n915), .B1(n84), .B2(n306), .ZN(n1107) );
  INV_X1 U436 ( .A(current_mask_in[1]), .ZN(n306) );
  OAI22_X1 U437 ( .A1(n77), .A2(n914), .B1(n84), .B2(n307), .ZN(n1106) );
  INV_X1 U438 ( .A(current_mask_in[2]), .ZN(n307) );
  OAI22_X1 U439 ( .A1(n77), .A2(n913), .B1(n85), .B2(n308), .ZN(n1105) );
  INV_X1 U440 ( .A(current_mask_in[3]), .ZN(n308) );
  OAI22_X1 U441 ( .A1(n78), .A2(n912), .B1(n85), .B2(n309), .ZN(n1104) );
  INV_X1 U442 ( .A(current_mask_in[4]), .ZN(n309) );
  OAI22_X1 U443 ( .A1(n78), .A2(n911), .B1(n85), .B2(n310), .ZN(n1103) );
  INV_X1 U444 ( .A(current_mask_in[5]), .ZN(n310) );
  OAI22_X1 U445 ( .A1(n78), .A2(n910), .B1(n85), .B2(n311), .ZN(n1102) );
  INV_X1 U446 ( .A(current_mask_in[6]), .ZN(n311) );
  OAI22_X1 U447 ( .A1(n78), .A2(n909), .B1(n85), .B2(n312), .ZN(n1101) );
  INV_X1 U448 ( .A(current_mask_in[7]), .ZN(n312) );
  OAI22_X1 U449 ( .A1(n78), .A2(n908), .B1(n85), .B2(n313), .ZN(n1100) );
  INV_X1 U450 ( .A(current_mask_in[8]), .ZN(n313) );
  OAI22_X1 U451 ( .A1(n78), .A2(n907), .B1(n85), .B2(n314), .ZN(n1099) );
  INV_X1 U452 ( .A(current_mask_in[9]), .ZN(n314) );
  OAI22_X1 U453 ( .A1(n78), .A2(n906), .B1(n85), .B2(n315), .ZN(n1098) );
  INV_X1 U454 ( .A(current_mask_in[10]), .ZN(n315) );
  OAI22_X1 U455 ( .A1(n78), .A2(n905), .B1(n85), .B2(n316), .ZN(n1097) );
  INV_X1 U456 ( .A(current_mask_in[11]), .ZN(n316) );
  OAI22_X1 U457 ( .A1(n78), .A2(n904), .B1(n85), .B2(n317), .ZN(n1096) );
  INV_X1 U458 ( .A(current_mask_in[12]), .ZN(n317) );
  OAI22_X1 U459 ( .A1(n78), .A2(n903), .B1(n85), .B2(n318), .ZN(n1095) );
  INV_X1 U460 ( .A(current_mask_in[13]), .ZN(n318) );
  OAI22_X1 U461 ( .A1(n78), .A2(n902), .B1(n85), .B2(n319), .ZN(n1094) );
  INV_X1 U462 ( .A(current_mask_in[14]), .ZN(n319) );
  OAI22_X1 U463 ( .A1(n78), .A2(n901), .B1(n86), .B2(n320), .ZN(n1093) );
  INV_X1 U464 ( .A(current_mask_in[15]), .ZN(n320) );
  OAI22_X1 U465 ( .A1(n79), .A2(n900), .B1(n86), .B2(n321), .ZN(n1092) );
  INV_X1 U466 ( .A(current_mask_in[16]), .ZN(n321) );
  OAI22_X1 U467 ( .A1(n79), .A2(n899), .B1(n86), .B2(n322), .ZN(n1091) );
  INV_X1 U468 ( .A(current_mask_in[17]), .ZN(n322) );
  OAI22_X1 U469 ( .A1(n79), .A2(n898), .B1(n86), .B2(n323), .ZN(n1090) );
  INV_X1 U470 ( .A(current_mask_in[18]), .ZN(n323) );
  OAI22_X1 U471 ( .A1(n79), .A2(n897), .B1(n86), .B2(n324), .ZN(n1089) );
  INV_X1 U472 ( .A(current_mask_in[19]), .ZN(n324) );
  OAI22_X1 U473 ( .A1(n79), .A2(n896), .B1(n86), .B2(n325), .ZN(n1088) );
  INV_X1 U474 ( .A(current_mask_in[20]), .ZN(n325) );
  OAI22_X1 U475 ( .A1(n79), .A2(n895), .B1(n86), .B2(n326), .ZN(n1087) );
  INV_X1 U476 ( .A(current_mask_in[21]), .ZN(n326) );
  OAI22_X1 U477 ( .A1(n79), .A2(n894), .B1(n86), .B2(n327), .ZN(n1086) );
  INV_X1 U478 ( .A(current_mask_in[22]), .ZN(n327) );
  OAI22_X1 U479 ( .A1(n79), .A2(n893), .B1(n86), .B2(n328), .ZN(n1085) );
  INV_X1 U480 ( .A(current_mask_in[23]), .ZN(n328) );
  OAI22_X1 U481 ( .A1(n79), .A2(n892), .B1(n86), .B2(n329), .ZN(n1084) );
  INV_X1 U482 ( .A(current_mask_in[24]), .ZN(n329) );
  OAI22_X1 U483 ( .A1(n79), .A2(n891), .B1(n86), .B2(n330), .ZN(n1083) );
  INV_X1 U484 ( .A(current_mask_in[25]), .ZN(n330) );
  OAI22_X1 U485 ( .A1(n79), .A2(n890), .B1(n86), .B2(n331), .ZN(n1082) );
  INV_X1 U486 ( .A(current_mask_in[26]), .ZN(n331) );
  OAI22_X1 U487 ( .A1(n79), .A2(n889), .B1(n87), .B2(n332), .ZN(n1081) );
  INV_X1 U488 ( .A(current_mask_in[27]), .ZN(n332) );
  OAI22_X1 U489 ( .A1(n79), .A2(n888), .B1(n87), .B2(n333), .ZN(n1080) );
  INV_X1 U490 ( .A(current_mask_in[28]), .ZN(n333) );
  OAI22_X1 U491 ( .A1(n82), .A2(n887), .B1(n87), .B2(n334), .ZN(n1079) );
  INV_X1 U492 ( .A(current_mask_in[29]), .ZN(n334) );
  OAI22_X1 U493 ( .A1(n81), .A2(n886), .B1(n87), .B2(n335), .ZN(n1078) );
  INV_X1 U494 ( .A(current_mask_in[30]), .ZN(n335) );
  OAI22_X1 U495 ( .A1(n80), .A2(n885), .B1(n87), .B2(n336), .ZN(n1077) );
  INV_X1 U496 ( .A(current_mask_in[31]), .ZN(n336) );
  OAI22_X1 U497 ( .A1(n78), .A2(n884), .B1(n87), .B2(n337), .ZN(n1076) );
  INV_X1 U498 ( .A(initial_mask_in[0]), .ZN(n337) );
  OAI22_X1 U499 ( .A1(n77), .A2(n883), .B1(n87), .B2(n338), .ZN(n1075) );
  INV_X1 U500 ( .A(initial_mask_in[1]), .ZN(n338) );
  OAI22_X1 U501 ( .A1(n79), .A2(n882), .B1(n87), .B2(n339), .ZN(n1074) );
  INV_X1 U502 ( .A(initial_mask_in[2]), .ZN(n339) );
  OAI22_X1 U503 ( .A1(n82), .A2(n881), .B1(n87), .B2(n340), .ZN(n1073) );
  INV_X1 U504 ( .A(initial_mask_in[3]), .ZN(n340) );
  OAI22_X1 U505 ( .A1(n81), .A2(n880), .B1(n87), .B2(n341), .ZN(n1072) );
  INV_X1 U506 ( .A(initial_mask_in[4]), .ZN(n341) );
  OAI22_X1 U507 ( .A1(n80), .A2(n879), .B1(n87), .B2(n342), .ZN(n1071) );
  INV_X1 U508 ( .A(initial_mask_in[5]), .ZN(n342) );
  OAI22_X1 U509 ( .A1(n81), .A2(n878), .B1(n87), .B2(n343), .ZN(n1070) );
  INV_X1 U510 ( .A(initial_mask_in[6]), .ZN(n343) );
  OAI22_X1 U511 ( .A1(n80), .A2(n877), .B1(n88), .B2(n344), .ZN(n1069) );
  INV_X1 U512 ( .A(initial_mask_in[7]), .ZN(n344) );
  OAI22_X1 U513 ( .A1(n77), .A2(n876), .B1(n88), .B2(n345), .ZN(n1068) );
  INV_X1 U514 ( .A(initial_mask_in[8]), .ZN(n345) );
  OAI22_X1 U515 ( .A1(n79), .A2(n875), .B1(n88), .B2(n346), .ZN(n1067) );
  INV_X1 U516 ( .A(initial_mask_in[9]), .ZN(n346) );
  OAI22_X1 U517 ( .A1(n81), .A2(n874), .B1(n88), .B2(n347), .ZN(n1066) );
  INV_X1 U518 ( .A(initial_mask_in[10]), .ZN(n347) );
  OAI22_X1 U519 ( .A1(n80), .A2(n873), .B1(n88), .B2(n348), .ZN(n1065) );
  INV_X1 U520 ( .A(initial_mask_in[11]), .ZN(n348) );
  OAI22_X1 U521 ( .A1(n77), .A2(n872), .B1(n88), .B2(n349), .ZN(n1064) );
  INV_X1 U522 ( .A(initial_mask_in[12]), .ZN(n349) );
  OAI22_X1 U523 ( .A1(n78), .A2(n871), .B1(n88), .B2(n350), .ZN(n1063) );
  INV_X1 U524 ( .A(initial_mask_in[13]), .ZN(n350) );
  OAI22_X1 U525 ( .A1(n77), .A2(n870), .B1(n88), .B2(n351), .ZN(n1062) );
  INV_X1 U526 ( .A(initial_mask_in[14]), .ZN(n351) );
  OAI22_X1 U527 ( .A1(n79), .A2(n869), .B1(n88), .B2(n352), .ZN(n1061) );
  INV_X1 U528 ( .A(initial_mask_in[15]), .ZN(n352) );
  OAI22_X1 U529 ( .A1(n81), .A2(n868), .B1(n88), .B2(n353), .ZN(n1060) );
  INV_X1 U530 ( .A(initial_mask_in[16]), .ZN(n353) );
  OAI22_X1 U531 ( .A1(n80), .A2(n867), .B1(n88), .B2(n354), .ZN(n1059) );
  INV_X1 U532 ( .A(initial_mask_in[17]), .ZN(n354) );
  OAI22_X1 U533 ( .A1(n79), .A2(n866), .B1(n89), .B2(n355), .ZN(n1058) );
  INV_X1 U534 ( .A(initial_mask_in[18]), .ZN(n355) );
  OAI22_X1 U535 ( .A1(n80), .A2(n865), .B1(n89), .B2(n356), .ZN(n1057) );
  INV_X1 U536 ( .A(initial_mask_in[19]), .ZN(n356) );
  OAI22_X1 U537 ( .A1(n80), .A2(n864), .B1(n89), .B2(n357), .ZN(n1056) );
  INV_X1 U538 ( .A(initial_mask_in[20]), .ZN(n357) );
  OAI22_X1 U539 ( .A1(n80), .A2(n863), .B1(n89), .B2(n358), .ZN(n1055) );
  INV_X1 U540 ( .A(initial_mask_in[21]), .ZN(n358) );
  OAI22_X1 U541 ( .A1(n80), .A2(n862), .B1(n89), .B2(n359), .ZN(n1054) );
  INV_X1 U542 ( .A(initial_mask_in[22]), .ZN(n359) );
  OAI22_X1 U543 ( .A1(n80), .A2(n861), .B1(n89), .B2(n360), .ZN(n1053) );
  INV_X1 U544 ( .A(initial_mask_in[23]), .ZN(n360) );
  OAI22_X1 U545 ( .A1(n80), .A2(n860), .B1(n89), .B2(n361), .ZN(n1052) );
  INV_X1 U546 ( .A(initial_mask_in[24]), .ZN(n361) );
  OAI22_X1 U547 ( .A1(n80), .A2(n859), .B1(n89), .B2(n362), .ZN(n1051) );
  INV_X1 U548 ( .A(initial_mask_in[25]), .ZN(n362) );
  OAI22_X1 U549 ( .A1(n80), .A2(n858), .B1(n89), .B2(n363), .ZN(n1050) );
  INV_X1 U550 ( .A(initial_mask_in[26]), .ZN(n363) );
  OAI22_X1 U551 ( .A1(n80), .A2(n857), .B1(n89), .B2(n364), .ZN(n1049) );
  INV_X1 U552 ( .A(initial_mask_in[27]), .ZN(n364) );
  OAI22_X1 U553 ( .A1(n80), .A2(n856), .B1(n89), .B2(n365), .ZN(n1048) );
  INV_X1 U554 ( .A(initial_mask_in[28]), .ZN(n365) );
  OAI22_X1 U555 ( .A1(n80), .A2(n855), .B1(n89), .B2(n366), .ZN(n1047) );
  INV_X1 U556 ( .A(initial_mask_in[29]), .ZN(n366) );
  OAI22_X1 U557 ( .A1(n80), .A2(n854), .B1(n90), .B2(n367), .ZN(n1046) );
  INV_X1 U558 ( .A(initial_mask_in[30]), .ZN(n367) );
  OAI22_X1 U559 ( .A1(n81), .A2(n853), .B1(n90), .B2(n368), .ZN(n1045) );
  INV_X1 U560 ( .A(initial_mask_in[31]), .ZN(n368) );
  OAI22_X1 U561 ( .A1(n81), .A2(n852), .B1(n90), .B2(n369), .ZN(n1044) );
  INV_X1 U562 ( .A(next_pc_in[0]), .ZN(n369) );
  OAI22_X1 U563 ( .A1(n81), .A2(n851), .B1(n90), .B2(n370), .ZN(n1043) );
  INV_X1 U564 ( .A(next_pc_in[1]), .ZN(n370) );
  OAI22_X1 U565 ( .A1(n81), .A2(n850), .B1(n90), .B2(n371), .ZN(n1042) );
  INV_X1 U566 ( .A(next_pc_in[2]), .ZN(n371) );
  OAI22_X1 U567 ( .A1(n81), .A2(n849), .B1(n90), .B2(n372), .ZN(n1041) );
  INV_X1 U568 ( .A(next_pc_in[3]), .ZN(n372) );
  OAI22_X1 U569 ( .A1(n81), .A2(n848), .B1(n90), .B2(n373), .ZN(n1040) );
  INV_X1 U570 ( .A(next_pc_in[4]), .ZN(n373) );
  OAI22_X1 U571 ( .A1(n81), .A2(n847), .B1(n90), .B2(n374), .ZN(n1039) );
  INV_X1 U572 ( .A(next_pc_in[5]), .ZN(n374) );
  OAI22_X1 U573 ( .A1(n81), .A2(n846), .B1(n90), .B2(n375), .ZN(n1038) );
  INV_X1 U574 ( .A(next_pc_in[6]), .ZN(n375) );
  OAI22_X1 U575 ( .A1(n81), .A2(n845), .B1(n90), .B2(n376), .ZN(n1037) );
  INV_X1 U576 ( .A(next_pc_in[7]), .ZN(n376) );
  OAI22_X1 U577 ( .A1(n81), .A2(n844), .B1(n90), .B2(n377), .ZN(n1036) );
  INV_X1 U578 ( .A(next_pc_in[8]), .ZN(n377) );
  OAI22_X1 U579 ( .A1(n81), .A2(n843), .B1(n90), .B2(n378), .ZN(n1035) );
  INV_X1 U580 ( .A(next_pc_in[9]), .ZN(n378) );
  OAI22_X1 U581 ( .A1(n81), .A2(n842), .B1(n91), .B2(n379), .ZN(n1034) );
  INV_X1 U582 ( .A(next_pc_in[10]), .ZN(n379) );
  OAI22_X1 U583 ( .A1(n81), .A2(n841), .B1(n91), .B2(n380), .ZN(n1033) );
  INV_X1 U584 ( .A(next_pc_in[11]), .ZN(n380) );
  OAI22_X1 U585 ( .A1(n80), .A2(n840), .B1(n91), .B2(n381), .ZN(n1032) );
  INV_X1 U586 ( .A(next_pc_in[12]), .ZN(n381) );
  OAI22_X1 U587 ( .A1(n77), .A2(n839), .B1(n91), .B2(n382), .ZN(n1031) );
  INV_X1 U588 ( .A(next_pc_in[13]), .ZN(n382) );
  OAI22_X1 U589 ( .A1(n79), .A2(n838), .B1(n91), .B2(n383), .ZN(n1030) );
  INV_X1 U590 ( .A(next_pc_in[14]), .ZN(n383) );
  OAI22_X1 U591 ( .A1(n82), .A2(n837), .B1(n91), .B2(n384), .ZN(n1029) );
  INV_X1 U592 ( .A(next_pc_in[15]), .ZN(n384) );
  OAI22_X1 U593 ( .A1(n81), .A2(n836), .B1(n91), .B2(n385), .ZN(n1028) );
  INV_X1 U594 ( .A(next_pc_in[16]), .ZN(n385) );
  OAI22_X1 U595 ( .A1(n80), .A2(n835), .B1(n91), .B2(n386), .ZN(n1027) );
  INV_X1 U596 ( .A(next_pc_in[17]), .ZN(n386) );
  OAI22_X1 U597 ( .A1(n77), .A2(n834), .B1(n91), .B2(n387), .ZN(n1026) );
  INV_X1 U598 ( .A(next_pc_in[18]), .ZN(n387) );
  OAI22_X1 U599 ( .A1(n79), .A2(n833), .B1(n91), .B2(n388), .ZN(n1025) );
  INV_X1 U600 ( .A(next_pc_in[19]), .ZN(n388) );
  OAI22_X1 U601 ( .A1(n82), .A2(n832), .B1(n91), .B2(n389), .ZN(n1024) );
  INV_X1 U602 ( .A(next_pc_in[20]), .ZN(n389) );
  OAI22_X1 U603 ( .A1(n81), .A2(n831), .B1(n91), .B2(n390), .ZN(n1023) );
  INV_X1 U604 ( .A(next_pc_in[21]), .ZN(n390) );
  OAI22_X1 U605 ( .A1(n80), .A2(n830), .B1(n92), .B2(n391), .ZN(n1022) );
  INV_X1 U606 ( .A(next_pc_in[22]), .ZN(n391) );
  OAI22_X1 U607 ( .A1(n82), .A2(n829), .B1(n92), .B2(n392), .ZN(n1021) );
  INV_X1 U608 ( .A(next_pc_in[23]), .ZN(n392) );
  OAI22_X1 U609 ( .A1(n82), .A2(n828), .B1(n92), .B2(n393), .ZN(n1020) );
  INV_X1 U610 ( .A(next_pc_in[24]), .ZN(n393) );
  OAI22_X1 U611 ( .A1(n82), .A2(n827), .B1(n92), .B2(n394), .ZN(n1019) );
  INV_X1 U612 ( .A(next_pc_in[25]), .ZN(n394) );
  OAI22_X1 U613 ( .A1(n82), .A2(n826), .B1(n92), .B2(n395), .ZN(n1018) );
  INV_X1 U614 ( .A(next_pc_in[26]), .ZN(n395) );
  OAI22_X1 U615 ( .A1(n82), .A2(n825), .B1(n92), .B2(n396), .ZN(n1017) );
  INV_X1 U616 ( .A(next_pc_in[27]), .ZN(n396) );
  OAI22_X1 U617 ( .A1(n82), .A2(n824), .B1(n92), .B2(n397), .ZN(n1016) );
  INV_X1 U618 ( .A(next_pc_in[28]), .ZN(n397) );
  OAI22_X1 U619 ( .A1(n82), .A2(n823), .B1(n92), .B2(n398), .ZN(n1015) );
  INV_X1 U620 ( .A(next_pc_in[29]), .ZN(n398) );
  OAI22_X1 U621 ( .A1(n82), .A2(n822), .B1(n92), .B2(n399), .ZN(n1014) );
  INV_X1 U622 ( .A(next_pc_in[30]), .ZN(n399) );
  OAI22_X1 U623 ( .A1(n82), .A2(n821), .B1(n92), .B2(n400), .ZN(n1013) );
  INV_X1 U624 ( .A(next_pc_in[31]), .ZN(n400) );
  OAI22_X1 U625 ( .A1(n82), .A2(n820), .B1(n92), .B2(n401), .ZN(n1012) );
  INV_X1 U626 ( .A(gprs_base_addr_in[0]), .ZN(n401) );
  OAI22_X1 U627 ( .A1(n82), .A2(n819), .B1(n92), .B2(n402), .ZN(n1011) );
  INV_X1 U628 ( .A(gprs_base_addr_in[1]), .ZN(n402) );
  OAI22_X1 U629 ( .A1(n81), .A2(n818), .B1(n93), .B2(n403), .ZN(n1010) );
  INV_X1 U630 ( .A(gprs_base_addr_in[2]), .ZN(n403) );
  OAI22_X1 U631 ( .A1(n82), .A2(n817), .B1(n93), .B2(n404), .ZN(n1009) );
  INV_X1 U632 ( .A(gprs_base_addr_in[3]), .ZN(n404) );
  OAI22_X1 U633 ( .A1(n82), .A2(n816), .B1(n93), .B2(n405), .ZN(n1008) );
  INV_X1 U634 ( .A(gprs_base_addr_in[4]), .ZN(n405) );
  OAI22_X1 U635 ( .A1(n80), .A2(n815), .B1(n93), .B2(n406), .ZN(n1007) );
  INV_X1 U636 ( .A(gprs_base_addr_in[5]), .ZN(n406) );
  OAI22_X1 U637 ( .A1(n78), .A2(n814), .B1(n93), .B2(n407), .ZN(n1006) );
  INV_X1 U638 ( .A(gprs_base_addr_in[6]), .ZN(n407) );
  OAI22_X1 U639 ( .A1(n82), .A2(n813), .B1(n93), .B2(n408), .ZN(n1005) );
  INV_X1 U640 ( .A(gprs_base_addr_in[7]), .ZN(n408) );
  OAI22_X1 U641 ( .A1(n79), .A2(n812), .B1(n93), .B2(n409), .ZN(n1004) );
  INV_X1 U642 ( .A(gprs_base_addr_in[8]), .ZN(n409) );
  OAI22_X1 U643 ( .A1(n77), .A2(n811), .B1(n93), .B2(n410), .ZN(n1003) );
  INV_X1 U644 ( .A(shmem_base_addr_in[0]), .ZN(n410) );
  OAI22_X1 U645 ( .A1(n78), .A2(n810), .B1(n93), .B2(n411), .ZN(n1002) );
  INV_X1 U646 ( .A(shmem_base_addr_in[1]), .ZN(n411) );
  OAI22_X1 U647 ( .A1(n77), .A2(n809), .B1(n93), .B2(n412), .ZN(n1001) );
  INV_X1 U648 ( .A(shmem_base_addr_in[2]), .ZN(n412) );
  OAI22_X1 U649 ( .A1(n77), .A2(n808), .B1(n83), .B2(n413), .ZN(n1000) );
  INV_X1 U650 ( .A(shmem_base_addr_in[3]), .ZN(n413) );
  NAND2_X1 U651 ( .A1(n181), .A2(n78), .ZN(n149) );
  NOR2_X1 U652 ( .A1(n304), .A2(n102), .ZN(n181) );
  OAI21_X1 U653 ( .B1(n182), .B2(n304), .A(n99), .ZN(n414) );
  INV_X1 U654 ( .A(en), .ZN(n304) );
  INV_X1 U655 ( .A(n302), .ZN(n182) );
  NAND2_X1 U656 ( .A1(warp_lane_id_in[1]), .A2(warp_lane_id_in[0]), .ZN(n302)
         );
  INV_X1 U657 ( .A(n257), .ZN(n187) );
  NOR3_X1 U658 ( .A1(warp_checker_state_machine[1]), .A2(
        warp_checker_state_machine[2]), .A3(n3), .ZN(n257) );
  INV_X1 U659 ( .A(n190), .ZN(n197) );
  NOR3_X1 U660 ( .A1(warp_checker_state_machine[0]), .A2(
        warp_checker_state_machine[1]), .A3(n8), .ZN(n190) );
  NOR2_X1 U661 ( .A1(n415), .A2(n416), .ZN(fence_id_mask[9]) );
  INV_X1 U662 ( .A(fence_regs_fence_en_in[9]), .ZN(n415) );
  NOR2_X1 U663 ( .A1(n417), .A2(n418), .ZN(fence_id_mask[8]) );
  INV_X1 U664 ( .A(fence_regs_fence_en_in[8]), .ZN(n417) );
  NOR2_X1 U665 ( .A1(n419), .A2(n420), .ZN(fence_id_mask[7]) );
  INV_X1 U666 ( .A(fence_regs_fence_en_in[7]), .ZN(n419) );
  NOR2_X1 U667 ( .A1(n421), .A2(n422), .ZN(fence_id_mask[6]) );
  INV_X1 U668 ( .A(fence_regs_fence_en_in[6]), .ZN(n421) );
  NOR2_X1 U669 ( .A1(n423), .A2(n424), .ZN(fence_id_mask[5]) );
  INV_X1 U670 ( .A(fence_regs_fence_en_in[5]), .ZN(n423) );
  NOR2_X1 U671 ( .A1(n425), .A2(n426), .ZN(fence_id_mask[4]) );
  INV_X1 U672 ( .A(fence_regs_fence_en_in[4]), .ZN(n425) );
  NOR2_X1 U673 ( .A1(n427), .A2(n428), .ZN(fence_id_mask[3]) );
  INV_X1 U674 ( .A(fence_regs_fence_en_in[3]), .ZN(n427) );
  NOR2_X1 U675 ( .A1(n429), .A2(n430), .ZN(fence_id_mask[31]) );
  INV_X1 U676 ( .A(fence_regs_fence_en_in[31]), .ZN(n429) );
  NOR2_X1 U677 ( .A1(n431), .A2(n432), .ZN(fence_id_mask[30]) );
  INV_X1 U678 ( .A(fence_regs_fence_en_in[30]), .ZN(n431) );
  NOR2_X1 U679 ( .A1(n433), .A2(n434), .ZN(fence_id_mask[2]) );
  INV_X1 U680 ( .A(fence_regs_fence_en_in[2]), .ZN(n433) );
  NOR2_X1 U681 ( .A1(n435), .A2(n436), .ZN(fence_id_mask[29]) );
  INV_X1 U682 ( .A(fence_regs_fence_en_in[29]), .ZN(n435) );
  NOR2_X1 U683 ( .A1(n437), .A2(n438), .ZN(fence_id_mask[28]) );
  INV_X1 U684 ( .A(fence_regs_fence_en_in[28]), .ZN(n437) );
  NOR2_X1 U685 ( .A1(n439), .A2(n440), .ZN(fence_id_mask[27]) );
  INV_X1 U686 ( .A(fence_regs_fence_en_in[27]), .ZN(n439) );
  NOR2_X1 U687 ( .A1(n441), .A2(n442), .ZN(fence_id_mask[26]) );
  INV_X1 U688 ( .A(fence_regs_fence_en_in[26]), .ZN(n441) );
  NOR2_X1 U689 ( .A1(n443), .A2(n444), .ZN(fence_id_mask[25]) );
  INV_X1 U690 ( .A(fence_regs_fence_en_in[25]), .ZN(n443) );
  NOR2_X1 U691 ( .A1(n445), .A2(n446), .ZN(fence_id_mask[24]) );
  INV_X1 U692 ( .A(fence_regs_fence_en_in[24]), .ZN(n445) );
  NOR2_X1 U693 ( .A1(n447), .A2(n448), .ZN(fence_id_mask[23]) );
  INV_X1 U694 ( .A(fence_regs_fence_en_in[23]), .ZN(n447) );
  NOR2_X1 U695 ( .A1(n449), .A2(n450), .ZN(fence_id_mask[22]) );
  INV_X1 U696 ( .A(fence_regs_fence_en_in[22]), .ZN(n449) );
  NOR2_X1 U697 ( .A1(n451), .A2(n452), .ZN(fence_id_mask[21]) );
  INV_X1 U698 ( .A(fence_regs_fence_en_in[21]), .ZN(n451) );
  NOR2_X1 U699 ( .A1(n453), .A2(n454), .ZN(fence_id_mask[20]) );
  INV_X1 U700 ( .A(fence_regs_fence_en_in[20]), .ZN(n453) );
  NOR2_X1 U701 ( .A1(n455), .A2(n456), .ZN(fence_id_mask[1]) );
  INV_X1 U702 ( .A(fence_regs_fence_en_in[1]), .ZN(n455) );
  NOR2_X1 U703 ( .A1(n457), .A2(n458), .ZN(fence_id_mask[19]) );
  INV_X1 U704 ( .A(fence_regs_fence_en_in[19]), .ZN(n457) );
  NOR2_X1 U705 ( .A1(n459), .A2(n460), .ZN(fence_id_mask[18]) );
  INV_X1 U706 ( .A(fence_regs_fence_en_in[18]), .ZN(n459) );
  NOR2_X1 U707 ( .A1(n461), .A2(n462), .ZN(fence_id_mask[17]) );
  INV_X1 U708 ( .A(fence_regs_fence_en_in[17]), .ZN(n461) );
  NOR2_X1 U709 ( .A1(n463), .A2(n464), .ZN(fence_id_mask[16]) );
  INV_X1 U710 ( .A(fence_regs_fence_en_in[16]), .ZN(n463) );
  NOR2_X1 U711 ( .A1(n465), .A2(n466), .ZN(fence_id_mask[15]) );
  INV_X1 U712 ( .A(fence_regs_fence_en_in[15]), .ZN(n465) );
  NOR2_X1 U713 ( .A1(n467), .A2(n468), .ZN(fence_id_mask[14]) );
  INV_X1 U714 ( .A(fence_regs_fence_en_in[14]), .ZN(n467) );
  NOR2_X1 U715 ( .A1(n469), .A2(n470), .ZN(fence_id_mask[13]) );
  INV_X1 U716 ( .A(fence_regs_fence_en_in[13]), .ZN(n469) );
  NOR2_X1 U717 ( .A1(n471), .A2(n472), .ZN(fence_id_mask[12]) );
  INV_X1 U718 ( .A(fence_regs_fence_en_in[12]), .ZN(n471) );
  NOR2_X1 U719 ( .A1(n473), .A2(n474), .ZN(fence_id_mask[11]) );
  INV_X1 U720 ( .A(fence_regs_fence_en_in[11]), .ZN(n473) );
  NOR2_X1 U721 ( .A1(n475), .A2(n476), .ZN(fence_id_mask[10]) );
  INV_X1 U722 ( .A(fence_regs_fence_en_in[10]), .ZN(n475) );
  NOR2_X1 U723 ( .A1(n477), .A2(n478), .ZN(fence_id_mask[0]) );
  INV_X1 U724 ( .A(fence_regs_fence_en_in[0]), .ZN(n477) );
  AOI21_X1 U725 ( .B1(n479), .B2(n480), .A(n416), .ZN(cta_id_mask_rev[9]) );
  NAND4_X1 U726 ( .A1(n481), .A2(n482), .A3(n483), .A4(n484), .ZN(n416) );
  XNOR2_X1 U727 ( .A(n137), .B(\fence_regs_cta_id_in[9><0] ), .ZN(n484) );
  XNOR2_X1 U728 ( .A(n139), .B(\fence_regs_cta_id_in[9><1] ), .ZN(n483) );
  XNOR2_X1 U729 ( .A(n141), .B(\fence_regs_cta_id_in[9><2] ), .ZN(n482) );
  XNOR2_X1 U730 ( .A(n143), .B(\fence_regs_cta_id_in[9><3] ), .ZN(n481) );
  AOI21_X1 U731 ( .B1(n479), .B2(n485), .A(n418), .ZN(cta_id_mask_rev[8]) );
  NAND4_X1 U732 ( .A1(n486), .A2(n487), .A3(n488), .A4(n489), .ZN(n418) );
  XNOR2_X1 U733 ( .A(n137), .B(\fence_regs_cta_id_in[8><0] ), .ZN(n489) );
  XNOR2_X1 U734 ( .A(n139), .B(\fence_regs_cta_id_in[8><1] ), .ZN(n488) );
  XNOR2_X1 U735 ( .A(n141), .B(\fence_regs_cta_id_in[8><2] ), .ZN(n487) );
  XNOR2_X1 U736 ( .A(n143), .B(\fence_regs_cta_id_in[8><3] ), .ZN(n486) );
  NOR2_X1 U737 ( .A1(n490), .A2(n420), .ZN(cta_id_mask_rev[7]) );
  NAND4_X1 U738 ( .A1(n491), .A2(n492), .A3(n493), .A4(n494), .ZN(n420) );
  XNOR2_X1 U739 ( .A(n137), .B(\fence_regs_cta_id_in[7><0] ), .ZN(n494) );
  XNOR2_X1 U740 ( .A(n139), .B(\fence_regs_cta_id_in[7><1] ), .ZN(n493) );
  XNOR2_X1 U741 ( .A(n141), .B(\fence_regs_cta_id_in[7><2] ), .ZN(n492) );
  XNOR2_X1 U742 ( .A(n143), .B(\fence_regs_cta_id_in[7><3] ), .ZN(n491) );
  NOR2_X1 U743 ( .A1(n495), .A2(n422), .ZN(cta_id_mask_rev[6]) );
  NAND4_X1 U744 ( .A1(n496), .A2(n497), .A3(n498), .A4(n499), .ZN(n422) );
  XNOR2_X1 U745 ( .A(n137), .B(\fence_regs_cta_id_in[6><0] ), .ZN(n499) );
  XNOR2_X1 U746 ( .A(n139), .B(\fence_regs_cta_id_in[6><1] ), .ZN(n498) );
  XNOR2_X1 U747 ( .A(n141), .B(\fence_regs_cta_id_in[6><2] ), .ZN(n497) );
  XNOR2_X1 U748 ( .A(n143), .B(\fence_regs_cta_id_in[6><3] ), .ZN(n496) );
  AOI21_X1 U749 ( .B1(n500), .B2(warps_per_block_in[2]), .A(n501), .ZN(n495)
         );
  NOR2_X1 U750 ( .A1(n502), .A2(n424), .ZN(cta_id_mask_rev[5]) );
  NAND4_X1 U751 ( .A1(n503), .A2(n504), .A3(n505), .A4(n506), .ZN(n424) );
  XNOR2_X1 U752 ( .A(n137), .B(\fence_regs_cta_id_in[5><0] ), .ZN(n506) );
  XNOR2_X1 U753 ( .A(n139), .B(\fence_regs_cta_id_in[5><1] ), .ZN(n505) );
  XNOR2_X1 U754 ( .A(n141), .B(\fence_regs_cta_id_in[5><2] ), .ZN(n504) );
  XNOR2_X1 U755 ( .A(n143), .B(\fence_regs_cta_id_in[5><3] ), .ZN(n503) );
  AOI21_X1 U756 ( .B1(warps_per_block_in[2]), .B2(warps_per_block_in[1]), .A(
        n501), .ZN(n502) );
  NOR2_X1 U757 ( .A1(n507), .A2(n426), .ZN(cta_id_mask_rev[4]) );
  NAND4_X1 U758 ( .A1(n508), .A2(n509), .A3(n510), .A4(n511), .ZN(n426) );
  XNOR2_X1 U759 ( .A(n137), .B(\fence_regs_cta_id_in[4><0] ), .ZN(n511) );
  XNOR2_X1 U760 ( .A(n139), .B(\fence_regs_cta_id_in[4><1] ), .ZN(n510) );
  XNOR2_X1 U761 ( .A(n141), .B(\fence_regs_cta_id_in[4><2] ), .ZN(n509) );
  XNOR2_X1 U762 ( .A(n143), .B(\fence_regs_cta_id_in[4><3] ), .ZN(n508) );
  AOI21_X1 U763 ( .B1(warps_per_block_in[2]), .B2(n512), .A(n501), .ZN(n507)
         );
  NOR2_X1 U764 ( .A1(n513), .A2(n428), .ZN(cta_id_mask_rev[3]) );
  NAND4_X1 U765 ( .A1(n514), .A2(n515), .A3(n516), .A4(n517), .ZN(n428) );
  XNOR2_X1 U766 ( .A(n137), .B(\fence_regs_cta_id_in[3><0] ), .ZN(n517) );
  XNOR2_X1 U767 ( .A(n139), .B(\fence_regs_cta_id_in[3><1] ), .ZN(n516) );
  XNOR2_X1 U768 ( .A(n141), .B(\fence_regs_cta_id_in[3><2] ), .ZN(n515) );
  XNOR2_X1 U769 ( .A(n143), .B(\fence_regs_cta_id_in[3><3] ), .ZN(n514) );
  NOR2_X1 U770 ( .A1(n518), .A2(n430), .ZN(cta_id_mask_rev[31]) );
  NAND4_X1 U771 ( .A1(n519), .A2(n520), .A3(n521), .A4(n522), .ZN(n430) );
  XNOR2_X1 U772 ( .A(n137), .B(\fence_regs_cta_id_in[31><0] ), .ZN(n522) );
  XNOR2_X1 U773 ( .A(n139), .B(\fence_regs_cta_id_in[31><1] ), .ZN(n521) );
  XNOR2_X1 U774 ( .A(n141), .B(\fence_regs_cta_id_in[31><2] ), .ZN(n520) );
  XNOR2_X1 U775 ( .A(n143), .B(\fence_regs_cta_id_in[31><3] ), .ZN(n519) );
  AOI21_X1 U776 ( .B1(n518), .B2(n523), .A(n432), .ZN(cta_id_mask_rev[30]) );
  NAND4_X1 U777 ( .A1(n524), .A2(n525), .A3(n526), .A4(n527), .ZN(n432) );
  XNOR2_X1 U778 ( .A(n137), .B(\fence_regs_cta_id_in[30><0] ), .ZN(n527) );
  XNOR2_X1 U779 ( .A(n139), .B(\fence_regs_cta_id_in[30><1] ), .ZN(n526) );
  XNOR2_X1 U780 ( .A(n141), .B(\fence_regs_cta_id_in[30><2] ), .ZN(n525) );
  XNOR2_X1 U781 ( .A(n143), .B(\fence_regs_cta_id_in[30><3] ), .ZN(n524) );
  NAND3_X1 U782 ( .A1(n528), .A2(warps_per_block_in[0]), .A3(n529), .ZN(n523)
         );
  AOI21_X1 U783 ( .B1(n530), .B2(n490), .A(n434), .ZN(cta_id_mask_rev[2]) );
  NAND4_X1 U784 ( .A1(n531), .A2(n532), .A3(n533), .A4(n534), .ZN(n434) );
  XNOR2_X1 U785 ( .A(n137), .B(\fence_regs_cta_id_in[2><0] ), .ZN(n534) );
  XNOR2_X1 U786 ( .A(n139), .B(\fence_regs_cta_id_in[2><1] ), .ZN(n533) );
  XNOR2_X1 U787 ( .A(n141), .B(\fence_regs_cta_id_in[2><2] ), .ZN(n532) );
  XNOR2_X1 U788 ( .A(n143), .B(\fence_regs_cta_id_in[2><3] ), .ZN(n531) );
  NOR2_X1 U789 ( .A1(n535), .A2(n436), .ZN(cta_id_mask_rev[29]) );
  NAND4_X1 U790 ( .A1(n536), .A2(n537), .A3(n538), .A4(n539), .ZN(n436) );
  XNOR2_X1 U791 ( .A(n137), .B(\fence_regs_cta_id_in[29><0] ), .ZN(n539) );
  XNOR2_X1 U792 ( .A(n139), .B(\fence_regs_cta_id_in[29><1] ), .ZN(n538) );
  XNOR2_X1 U793 ( .A(n141), .B(\fence_regs_cta_id_in[29><2] ), .ZN(n537) );
  XNOR2_X1 U794 ( .A(n143), .B(\fence_regs_cta_id_in[29><3] ), .ZN(n536) );
  AOI21_X1 U795 ( .B1(n529), .B2(n528), .A(n540), .ZN(n535) );
  NOR2_X1 U796 ( .A1(n541), .A2(n438), .ZN(cta_id_mask_rev[28]) );
  NAND4_X1 U797 ( .A1(n542), .A2(n543), .A3(n544), .A4(n545), .ZN(n438) );
  XNOR2_X1 U798 ( .A(n137), .B(\fence_regs_cta_id_in[28><0] ), .ZN(n545) );
  XNOR2_X1 U799 ( .A(n139), .B(\fence_regs_cta_id_in[28><1] ), .ZN(n544) );
  XNOR2_X1 U800 ( .A(n141), .B(\fence_regs_cta_id_in[28><2] ), .ZN(n543) );
  XNOR2_X1 U801 ( .A(n143), .B(\fence_regs_cta_id_in[28><3] ), .ZN(n542) );
  AOI21_X1 U802 ( .B1(n546), .B2(n529), .A(n540), .ZN(n541) );
  NOR2_X1 U803 ( .A1(n547), .A2(n440), .ZN(cta_id_mask_rev[27]) );
  NAND4_X1 U804 ( .A1(n548), .A2(n549), .A3(n550), .A4(n551), .ZN(n440) );
  XNOR2_X1 U805 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[27><0] ), .ZN(
        n551) );
  XNOR2_X1 U806 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[27><1] ), .ZN(
        n550) );
  XNOR2_X1 U807 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[27><2] ), .ZN(
        n549) );
  XNOR2_X1 U808 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[27><3] ), .ZN(
        n548) );
  AOI21_X1 U809 ( .B1(n518), .B2(n552), .A(n442), .ZN(cta_id_mask_rev[26]) );
  NAND4_X1 U810 ( .A1(n553), .A2(n554), .A3(n555), .A4(n556), .ZN(n442) );
  XNOR2_X1 U811 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[26><0] ), .ZN(
        n556) );
  XNOR2_X1 U812 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[26><1] ), .ZN(
        n555) );
  XNOR2_X1 U813 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[26><2] ), .ZN(
        n554) );
  XNOR2_X1 U814 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[26><3] ), .ZN(
        n553) );
  NAND3_X1 U815 ( .A1(warps_per_block_in[3]), .A2(n557), .A3(
        warps_per_block_in[4]), .ZN(n552) );
  INV_X1 U816 ( .A(n540), .ZN(n518) );
  AOI21_X1 U817 ( .B1(n547), .B2(n558), .A(n444), .ZN(cta_id_mask_rev[25]) );
  NAND4_X1 U818 ( .A1(n559), .A2(n560), .A3(n561), .A4(n562), .ZN(n444) );
  XNOR2_X1 U819 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[25><0] ), .ZN(
        n562) );
  XNOR2_X1 U820 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[25><1] ), .ZN(
        n561) );
  XNOR2_X1 U821 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[25><2] ), .ZN(
        n560) );
  XNOR2_X1 U822 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[25><3] ), .ZN(
        n559) );
  NAND2_X1 U823 ( .A1(n528), .A2(warps_per_block_in[4]), .ZN(n558) );
  AOI21_X1 U824 ( .B1(n547), .B2(n563), .A(n446), .ZN(cta_id_mask_rev[24]) );
  NAND4_X1 U825 ( .A1(n564), .A2(n565), .A3(n566), .A4(n567), .ZN(n446) );
  XNOR2_X1 U826 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[24><0] ), .ZN(
        n567) );
  XNOR2_X1 U827 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[24><1] ), .ZN(
        n566) );
  XNOR2_X1 U828 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[24><2] ), .ZN(
        n565) );
  XNOR2_X1 U829 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[24><3] ), .ZN(
        n564) );
  NAND2_X1 U830 ( .A1(n546), .A2(warps_per_block_in[4]), .ZN(n563) );
  AOI21_X1 U831 ( .B1(warps_per_block_in[3]), .B2(n529), .A(n540), .ZN(n547)
         );
  NOR2_X1 U832 ( .A1(n568), .A2(n448), .ZN(cta_id_mask_rev[23]) );
  NAND4_X1 U833 ( .A1(n569), .A2(n570), .A3(n571), .A4(n572), .ZN(n448) );
  XNOR2_X1 U834 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[23><0] ), .ZN(
        n572) );
  XNOR2_X1 U835 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[23><1] ), .ZN(
        n571) );
  XNOR2_X1 U836 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[23><2] ), .ZN(
        n570) );
  XNOR2_X1 U837 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[23><3] ), .ZN(
        n569) );
  AOI21_X1 U838 ( .B1(n568), .B2(n573), .A(n450), .ZN(cta_id_mask_rev[22]) );
  NAND4_X1 U839 ( .A1(n574), .A2(n575), .A3(n576), .A4(n577), .ZN(n450) );
  XNOR2_X1 U840 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[22><0] ), .ZN(
        n577) );
  XNOR2_X1 U841 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[22><1] ), .ZN(
        n576) );
  XNOR2_X1 U842 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[22><2] ), .ZN(
        n575) );
  XNOR2_X1 U843 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[22><3] ), .ZN(
        n574) );
  NAND2_X1 U844 ( .A1(n529), .A2(n500), .ZN(n573) );
  AOI21_X1 U845 ( .B1(n568), .B2(n578), .A(n452), .ZN(cta_id_mask_rev[21]) );
  NAND4_X1 U846 ( .A1(n579), .A2(n580), .A3(n581), .A4(n582), .ZN(n452) );
  XNOR2_X1 U847 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[21><0] ), .ZN(
        n582) );
  XNOR2_X1 U848 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[21><1] ), .ZN(
        n581) );
  XNOR2_X1 U849 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[21><2] ), .ZN(
        n580) );
  XNOR2_X1 U850 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[21><3] ), .ZN(
        n579) );
  NAND2_X1 U851 ( .A1(n529), .A2(warps_per_block_in[1]), .ZN(n578) );
  AOI21_X1 U852 ( .B1(n568), .B2(n583), .A(n454), .ZN(cta_id_mask_rev[20]) );
  NAND4_X1 U853 ( .A1(n584), .A2(n585), .A3(n586), .A4(n587), .ZN(n454) );
  XNOR2_X1 U854 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[20><0] ), .ZN(
        n587) );
  XNOR2_X1 U855 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[20><1] ), .ZN(
        n586) );
  XNOR2_X1 U856 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[20><2] ), .ZN(
        n585) );
  XNOR2_X1 U857 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[20><3] ), .ZN(
        n584) );
  NAND2_X1 U858 ( .A1(n529), .A2(n512), .ZN(n583) );
  INV_X1 U859 ( .A(n588), .ZN(n529) );
  AOI21_X1 U860 ( .B1(n513), .B2(n589), .A(n456), .ZN(cta_id_mask_rev[1]) );
  NAND4_X1 U861 ( .A1(n590), .A2(n591), .A3(n592), .A4(n593), .ZN(n456) );
  XNOR2_X1 U862 ( .A(n137), .B(\fence_regs_cta_id_in[1><0] ), .ZN(n593) );
  XNOR2_X1 U863 ( .A(n139), .B(\fence_regs_cta_id_in[1><1] ), .ZN(n592) );
  XNOR2_X1 U864 ( .A(n141), .B(\fence_regs_cta_id_in[1><2] ), .ZN(n591) );
  XNOR2_X1 U865 ( .A(n143), .B(\fence_regs_cta_id_in[1><3] ), .ZN(n590) );
  INV_X1 U866 ( .A(warps_per_block_in[1]), .ZN(n589) );
  NOR2_X1 U867 ( .A1(n594), .A2(n458), .ZN(cta_id_mask_rev[19]) );
  NAND4_X1 U868 ( .A1(n595), .A2(n596), .A3(n597), .A4(n598), .ZN(n458) );
  XNOR2_X1 U869 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[19><0] ), .ZN(
        n598) );
  XNOR2_X1 U870 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[19><1] ), .ZN(
        n597) );
  XNOR2_X1 U871 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[19><2] ), .ZN(
        n596) );
  XNOR2_X1 U872 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[19><3] ), .ZN(
        n595) );
  INV_X1 U873 ( .A(n599), .ZN(n594) );
  AOI21_X1 U874 ( .B1(n568), .B2(n600), .A(n460), .ZN(cta_id_mask_rev[18]) );
  NAND4_X1 U875 ( .A1(n601), .A2(n602), .A3(n603), .A4(n604), .ZN(n460) );
  XNOR2_X1 U876 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[18><0] ), .ZN(
        n604) );
  XNOR2_X1 U877 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[18><1] ), .ZN(
        n603) );
  XNOR2_X1 U878 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[18><2] ), .ZN(
        n602) );
  XNOR2_X1 U879 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[18><3] ), .ZN(
        n601) );
  NAND2_X1 U880 ( .A1(warps_per_block_in[4]), .A2(n557), .ZN(n600) );
  NOR2_X1 U881 ( .A1(n605), .A2(n462), .ZN(cta_id_mask_rev[17]) );
  NAND4_X1 U882 ( .A1(n606), .A2(n607), .A3(n608), .A4(n609), .ZN(n462) );
  XNOR2_X1 U883 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[17><0] ), .ZN(
        n609) );
  XNOR2_X1 U884 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[17><1] ), .ZN(
        n608) );
  XNOR2_X1 U885 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[17><2] ), .ZN(
        n607) );
  XNOR2_X1 U886 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[17><3] ), .ZN(
        n606) );
  AOI21_X1 U887 ( .B1(warps_per_block_in[4]), .B2(warps_per_block_in[1]), .A(
        n599), .ZN(n605) );
  NOR2_X1 U888 ( .A1(n610), .A2(n464), .ZN(cta_id_mask_rev[16]) );
  NAND4_X1 U889 ( .A1(n611), .A2(n612), .A3(n613), .A4(n614), .ZN(n464) );
  XNOR2_X1 U890 ( .A(n137), .B(\fence_regs_cta_id_in[16><0] ), .ZN(n614) );
  XNOR2_X1 U891 ( .A(n139), .B(\fence_regs_cta_id_in[16><1] ), .ZN(n613) );
  XNOR2_X1 U892 ( .A(n141), .B(\fence_regs_cta_id_in[16><2] ), .ZN(n612) );
  XNOR2_X1 U893 ( .A(n143), .B(\fence_regs_cta_id_in[16><3] ), .ZN(n611) );
  AOI21_X1 U894 ( .B1(warps_per_block_in[4]), .B2(n512), .A(n599), .ZN(n610)
         );
  NAND2_X1 U895 ( .A1(n568), .A2(n588), .ZN(n599) );
  NAND2_X1 U896 ( .A1(warps_per_block_in[4]), .A2(warps_per_block_in[2]), .ZN(
        n588) );
  AOI21_X1 U897 ( .B1(warps_per_block_in[3]), .B2(warps_per_block_in[4]), .A(
        n540), .ZN(n568) );
  NOR2_X1 U898 ( .A1(n615), .A2(n466), .ZN(cta_id_mask_rev[15]) );
  NAND4_X1 U899 ( .A1(n616), .A2(n617), .A3(n618), .A4(n619), .ZN(n466) );
  XNOR2_X1 U900 ( .A(n137), .B(\fence_regs_cta_id_in[15><0] ), .ZN(n619) );
  XNOR2_X1 U901 ( .A(n139), .B(\fence_regs_cta_id_in[15><1] ), .ZN(n618) );
  XNOR2_X1 U902 ( .A(n141), .B(\fence_regs_cta_id_in[15><2] ), .ZN(n617) );
  XNOR2_X1 U903 ( .A(n143), .B(\fence_regs_cta_id_in[15><3] ), .ZN(n616) );
  AOI21_X1 U904 ( .B1(n615), .B2(n620), .A(n468), .ZN(cta_id_mask_rev[14]) );
  NAND4_X1 U905 ( .A1(n621), .A2(n622), .A3(n623), .A4(n624), .ZN(n468) );
  XNOR2_X1 U906 ( .A(n137), .B(\fence_regs_cta_id_in[14><0] ), .ZN(n624) );
  XNOR2_X1 U907 ( .A(n139), .B(\fence_regs_cta_id_in[14><1] ), .ZN(n623) );
  XNOR2_X1 U908 ( .A(n141), .B(\fence_regs_cta_id_in[14><2] ), .ZN(n622) );
  XNOR2_X1 U909 ( .A(n143), .B(\fence_regs_cta_id_in[14><3] ), .ZN(n621) );
  NAND3_X1 U910 ( .A1(warps_per_block_in[0]), .A2(warps_per_block_in[2]), .A3(
        n528), .ZN(n620) );
  AOI21_X1 U911 ( .B1(n615), .B2(n625), .A(n470), .ZN(cta_id_mask_rev[13]) );
  NAND4_X1 U912 ( .A1(n626), .A2(n627), .A3(n628), .A4(n629), .ZN(n470) );
  XNOR2_X1 U913 ( .A(n137), .B(\fence_regs_cta_id_in[13><0] ), .ZN(n629) );
  XNOR2_X1 U914 ( .A(n139), .B(\fence_regs_cta_id_in[13><1] ), .ZN(n628) );
  XNOR2_X1 U915 ( .A(n141), .B(\fence_regs_cta_id_in[13><2] ), .ZN(n627) );
  XNOR2_X1 U916 ( .A(n143), .B(\fence_regs_cta_id_in[13><3] ), .ZN(n626) );
  NAND2_X1 U917 ( .A1(n528), .A2(warps_per_block_in[2]), .ZN(n625) );
  INV_X1 U918 ( .A(n480), .ZN(n528) );
  NAND2_X1 U919 ( .A1(warps_per_block_in[3]), .A2(warps_per_block_in[1]), .ZN(
        n480) );
  AOI21_X1 U920 ( .B1(n615), .B2(n630), .A(n472), .ZN(cta_id_mask_rev[12]) );
  NAND4_X1 U921 ( .A1(n631), .A2(n632), .A3(n633), .A4(n634), .ZN(n472) );
  XNOR2_X1 U922 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[12><0] ), .ZN(
        n634) );
  XNOR2_X1 U923 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[12><1] ), .ZN(
        n633) );
  XNOR2_X1 U924 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[12><2] ), .ZN(
        n632) );
  XNOR2_X1 U925 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[12><3] ), .ZN(
        n631) );
  NAND2_X1 U926 ( .A1(n546), .A2(warps_per_block_in[2]), .ZN(n630) );
  INV_X1 U927 ( .A(n485), .ZN(n546) );
  NAND2_X1 U928 ( .A1(warps_per_block_in[3]), .A2(n512), .ZN(n485) );
  INV_X1 U929 ( .A(n635), .ZN(n512) );
  NOR2_X1 U930 ( .A1(n479), .A2(n474), .ZN(cta_id_mask_rev[11]) );
  NAND4_X1 U931 ( .A1(n636), .A2(n637), .A3(n638), .A4(n639), .ZN(n474) );
  XNOR2_X1 U932 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[11><0] ), .ZN(
        n639) );
  XNOR2_X1 U933 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[11><1] ), .ZN(
        n638) );
  XNOR2_X1 U934 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[11><2] ), .ZN(
        n637) );
  XNOR2_X1 U935 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[11><3] ), .ZN(
        n636) );
  AOI21_X1 U936 ( .B1(warps_per_block_in[3]), .B2(warps_per_block_in[2]), .A(
        n640), .ZN(n479) );
  AOI21_X1 U937 ( .B1(n615), .B2(n641), .A(n476), .ZN(cta_id_mask_rev[10]) );
  NAND4_X1 U938 ( .A1(n642), .A2(n643), .A3(n644), .A4(n645), .ZN(n476) );
  XNOR2_X1 U939 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[10><0] ), .ZN(
        n645) );
  XNOR2_X1 U940 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[10><1] ), .ZN(
        n644) );
  XNOR2_X1 U941 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[10><2] ), .ZN(
        n643) );
  XNOR2_X1 U942 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[10><3] ), .ZN(
        n642) );
  NAND2_X1 U943 ( .A1(warps_per_block_in[3]), .A2(n557), .ZN(n641) );
  INV_X1 U944 ( .A(n530), .ZN(n557) );
  NOR2_X1 U945 ( .A1(warps_per_block_in[2]), .A2(n500), .ZN(n530) );
  AND2_X1 U946 ( .A1(warps_per_block_in[0]), .A2(warps_per_block_in[1]), .ZN(
        n500) );
  AOI21_X1 U947 ( .B1(n635), .B2(n513), .A(n478), .ZN(cta_id_mask_rev[0]) );
  NAND4_X1 U948 ( .A1(n646), .A2(n647), .A3(n648), .A4(n649), .ZN(n478) );
  XNOR2_X1 U949 ( .A(n137), .B(\fence_regs_cta_id_in[0><0] ), .ZN(n649) );
  XNOR2_X1 U950 ( .A(n139), .B(\fence_regs_cta_id_in[0><1] ), .ZN(n648) );
  XNOR2_X1 U951 ( .A(n141), .B(\fence_regs_cta_id_in[0><2] ), .ZN(n647) );
  XNOR2_X1 U952 ( .A(n143), .B(\fence_regs_cta_id_in[0><3] ), .ZN(n646) );
  NOR2_X1 U953 ( .A1(n501), .A2(warps_per_block_in[2]), .ZN(n513) );
  INV_X1 U954 ( .A(n490), .ZN(n501) );
  NOR2_X1 U955 ( .A1(n640), .A2(warps_per_block_in[3]), .ZN(n490) );
  INV_X1 U956 ( .A(n615), .ZN(n640) );
  NOR2_X1 U957 ( .A1(n540), .A2(warps_per_block_in[4]), .ZN(n615) );
  NAND4_X1 U958 ( .A1(n142), .A2(n144), .A3(n140), .A4(n650), .ZN(n540) );
  NOR2_X1 U959 ( .A1(cta_id_in[0]), .A2(N1190), .ZN(n650) );
  NOR2_X1 U960 ( .A1(warps_per_block_in[1]), .A2(warps_per_block_in[0]), .ZN(
        n635) );
endmodule






module warp_generator_SHMEM_ADDR_SIZE14_DW01_inc_1 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(carry[11]), .B(A[11]), .Z(SUM[11]) );
  INV_X1 U2 ( .A(A[0]), .ZN(SUM[0]) );
endmodule


module warp_generator_SHMEM_ADDR_SIZE14_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  OR2_X1 U2 ( .A1(B[3]), .A2(A[3]), .ZN(n1) );
  INV_X1 U3 ( .A(n19), .ZN(n7) );
  INV_X1 U4 ( .A(n41), .ZN(n5) );
  INV_X1 U5 ( .A(n28), .ZN(n10) );
  INV_X1 U6 ( .A(n44), .ZN(n8) );
  INV_X1 U7 ( .A(n35), .ZN(n11) );
  INV_X1 U8 ( .A(n30), .ZN(n9) );
  INV_X1 U9 ( .A(A[2]), .ZN(n12) );
  INV_X1 U10 ( .A(n16), .ZN(n6) );
  AND2_X1 U11 ( .A1(n36), .A2(n1), .ZN(SUM[3]) );
  BUF_X1 U12 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  XOR2_X1 U14 ( .A(n13), .B(n14), .Z(SUM[9]) );
  NAND2_X1 U15 ( .A1(n15), .A2(n6), .ZN(n13) );
  XOR2_X1 U16 ( .A(n17), .B(n18), .Z(SUM[8]) );
  NOR2_X1 U17 ( .A1(n19), .A2(n20), .ZN(n18) );
  XNOR2_X1 U18 ( .A(n21), .B(n22), .ZN(SUM[7]) );
  AND2_X1 U19 ( .A1(n23), .A2(n8), .ZN(n22) );
  AOI21_X1 U20 ( .B1(n24), .B2(n25), .A(n9), .ZN(n21) );
  XNOR2_X1 U21 ( .A(n26), .B(n24), .ZN(SUM[6]) );
  OAI21_X1 U22 ( .B1(n27), .B2(n28), .A(n29), .ZN(n24) );
  NAND2_X1 U23 ( .A1(n25), .A2(n30), .ZN(n26) );
  XNOR2_X1 U24 ( .A(n27), .B(n31), .ZN(SUM[5]) );
  AND2_X1 U25 ( .A1(n29), .A2(n10), .ZN(n31) );
  NOR2_X1 U26 ( .A1(n32), .A2(n11), .ZN(n27) );
  XNOR2_X1 U27 ( .A(n36), .B(n33), .ZN(SUM[4]) );
  NOR2_X1 U28 ( .A1(n34), .A2(n11), .ZN(n33) );
  INV_X1 U29 ( .A(n12), .ZN(SUM[2]) );
  XOR2_X1 U30 ( .A(n37), .B(n38), .Z(SUM[11]) );
  AOI21_X1 U31 ( .B1(n39), .B2(n5), .A(n40), .ZN(n38) );
  XNOR2_X1 U32 ( .A(B[11]), .B(A[11]), .ZN(n37) );
  XOR2_X1 U33 ( .A(n39), .B(n42), .Z(SUM[10]) );
  NOR2_X1 U34 ( .A1(n41), .A2(n40), .ZN(n42) );
  AND2_X1 U35 ( .A1(B[10]), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U36 ( .A1(B[10]), .A2(A[10]), .ZN(n41) );
  OAI21_X1 U37 ( .B1(n16), .B2(n14), .A(n15), .ZN(n39) );
  NAND2_X1 U38 ( .A1(B[9]), .A2(A[9]), .ZN(n15) );
  AOI21_X1 U39 ( .B1(n7), .B2(n17), .A(n20), .ZN(n14) );
  AND2_X1 U40 ( .A1(B[8]), .A2(A[8]), .ZN(n20) );
  OAI211_X1 U41 ( .C1(n43), .C2(n44), .A(n23), .B(n45), .ZN(n17) );
  NAND4_X1 U42 ( .A1(n32), .A2(n10), .A3(n25), .A4(n8), .ZN(n45) );
  NOR2_X1 U43 ( .A1(n36), .A2(n34), .ZN(n32) );
  NOR2_X1 U44 ( .A1(B[4]), .A2(A[4]), .ZN(n34) );
  NAND2_X1 U45 ( .A1(B[3]), .A2(A[3]), .ZN(n36) );
  NAND2_X1 U46 ( .A1(B[7]), .A2(A[7]), .ZN(n23) );
  NOR2_X1 U47 ( .A1(B[7]), .A2(A[7]), .ZN(n44) );
  AOI21_X1 U48 ( .B1(n25), .B2(n46), .A(n9), .ZN(n43) );
  NAND2_X1 U49 ( .A1(B[6]), .A2(A[6]), .ZN(n30) );
  OAI21_X1 U50 ( .B1(n28), .B2(n35), .A(n29), .ZN(n46) );
  NAND2_X1 U51 ( .A1(B[5]), .A2(A[5]), .ZN(n29) );
  NAND2_X1 U52 ( .A1(B[4]), .A2(A[4]), .ZN(n35) );
  NOR2_X1 U53 ( .A1(B[5]), .A2(A[5]), .ZN(n28) );
  OR2_X1 U54 ( .A1(B[6]), .A2(A[6]), .ZN(n25) );
  NOR2_X1 U55 ( .A1(B[8]), .A2(A[8]), .ZN(n19) );
  NOR2_X1 U56 ( .A1(B[9]), .A2(A[9]), .ZN(n16) );
endmodule


module warp_generator_SHMEM_ADDR_SIZE14_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [3:0] A;
  input [13:0] B;
  output [17:0] PRODUCT;
  input TC;
  wire   \ab[3><13] , \ab[3><12] , \ab[3><11] , \ab[3><10] , \ab[3><9] ,
         \ab[3><8] , \ab[3><7] , \ab[3><6] , \ab[3><5] , \ab[3><4] ,
         \ab[3><3] , \ab[3><2] , \ab[3><1] , \ab[3><0] , \ab[2><13] ,
         \ab[2><12] , \ab[2><11] , \ab[2><10] , \ab[2><9] , \ab[2><8] ,
         \ab[2><7] , \ab[2><6] , \ab[2><5] , \ab[2><4] , \ab[2><3] ,
         \ab[2><2] , \ab[2><1] , \ab[2><0] , \ab[1><13] , \ab[1><12] ,
         \ab[1><11] , \ab[1><10] , \ab[1><9] , \ab[1><8] , \ab[1><7] ,
         \ab[1><6] , \ab[1><5] , \ab[1><4] , \ab[1><3] , \ab[1><2] ,
         \ab[1><1] , \ab[1><0] , \ab[0><13] , \ab[0><12] , \ab[0><11] ,
         \ab[0><10] , \ab[0><9] , \ab[0><8] , \ab[0><7] , \ab[0><6] ,
         \ab[0><5] , \ab[0><4] , \ab[0><3] , \ab[0><2] , \ab[0><1] ,
         \CARRYB[3><12] , \CARRYB[3><11] , \CARRYB[3><10] , \CARRYB[3><9] ,
         \CARRYB[3><8] , \CARRYB[3><7] , \CARRYB[3><6] , \CARRYB[3><5] ,
         \CARRYB[3><4] , \CARRYB[3><3] , \CARRYB[3><2] , \CARRYB[3><1] ,
         \CARRYB[3><0] , \CARRYB[2><12] , \CARRYB[2><11] , \CARRYB[2><10] ,
         \CARRYB[2><9] , \CARRYB[2><8] , \CARRYB[2><7] , \CARRYB[2><6] ,
         \CARRYB[2><5] , \CARRYB[2><4] , \CARRYB[2><3] , \CARRYB[2><2] ,
         \CARRYB[2><1] , \CARRYB[2><0] , \SUMB[3><12] , \SUMB[3><11] ,
         \SUMB[3><10] , \SUMB[3><9] , \SUMB[3><8] , \SUMB[3><7] , \SUMB[3><6] ,
         \SUMB[3><5] , \SUMB[3><4] , \SUMB[3><3] , \SUMB[3><2] , \SUMB[3><1] ,
         \SUMB[3><0] , \SUMB[2><12] , \SUMB[2><11] , \SUMB[2><10] ,
         \SUMB[2><9] , \SUMB[2><8] , \SUMB[2><7] , \SUMB[2><6] , \SUMB[2><5] ,
         \SUMB[2><4] , \SUMB[2><3] , \SUMB[2><2] , \SUMB[2><1] , \A1[0] , n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  FA_X1 S4_0 ( .A(\ab[3><0] ), .B(\CARRYB[2><0] ), .CI(\SUMB[2><1] ), .CO(
        \CARRYB[3><0] ), .S(\SUMB[3><0] ) );
  FA_X1 S4_1 ( .A(\ab[3><1] ), .B(\CARRYB[2><1] ), .CI(\SUMB[2><2] ), .CO(
        \CARRYB[3><1] ), .S(\SUMB[3><1] ) );
  FA_X1 S4_2 ( .A(\ab[3><2] ), .B(\CARRYB[2><2] ), .CI(\SUMB[2><3] ), .CO(
        \CARRYB[3><2] ), .S(\SUMB[3><2] ) );
  FA_X1 S4_3 ( .A(\ab[3><3] ), .B(\CARRYB[2><3] ), .CI(\SUMB[2><4] ), .CO(
        \CARRYB[3><3] ), .S(\SUMB[3><3] ) );
  FA_X1 S4_4 ( .A(\ab[3><4] ), .B(\CARRYB[2><4] ), .CI(\SUMB[2><5] ), .CO(
        \CARRYB[3><4] ), .S(\SUMB[3><4] ) );
  FA_X1 S4_5 ( .A(\ab[3><5] ), .B(\CARRYB[2><5] ), .CI(\SUMB[2><6] ), .CO(
        \CARRYB[3><5] ), .S(\SUMB[3><5] ) );
  FA_X1 S4_6 ( .A(\ab[3><6] ), .B(\CARRYB[2><6] ), .CI(\SUMB[2><7] ), .CO(
        \CARRYB[3><6] ), .S(\SUMB[3><6] ) );
  FA_X1 S4_7 ( .A(\ab[3><7] ), .B(\CARRYB[2><7] ), .CI(\SUMB[2><8] ), .CO(
        \CARRYB[3><7] ), .S(\SUMB[3><7] ) );
  FA_X1 S4_8 ( .A(\ab[3><8] ), .B(\CARRYB[2><8] ), .CI(\SUMB[2><9] ), .CO(
        \CARRYB[3><8] ), .S(\SUMB[3><8] ) );
  FA_X1 S4_9 ( .A(\ab[3><9] ), .B(\CARRYB[2><9] ), .CI(\SUMB[2><10] ), .CO(
        \CARRYB[3><9] ), .S(\SUMB[3><9] ) );
  FA_X1 S4_10 ( .A(\ab[3><10] ), .B(\CARRYB[2><10] ), .CI(\SUMB[2><11] ), .CO(
        \CARRYB[3><10] ), .S(\SUMB[3><10] ) );
  FA_X1 S4_11 ( .A(\ab[3><11] ), .B(\CARRYB[2><11] ), .CI(\SUMB[2><12] ), .CO(
        \CARRYB[3><11] ), .S(\SUMB[3><11] ) );
  FA_X1 S5_12 ( .A(\ab[3><12] ), .B(\CARRYB[2><12] ), .CI(\ab[2><13] ), .CO(
        \CARRYB[3><12] ), .S(\SUMB[3><12] ) );
  FA_X1 S1_2_0 ( .A(\ab[2><0] ), .B(n20), .CI(n34), .CO(\CARRYB[2><0] ), .S(
        \A1[0] ) );
  FA_X1 S2_2_1 ( .A(\ab[2><1] ), .B(n19), .CI(n33), .CO(\CARRYB[2><1] ), .S(
        \SUMB[2><1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2><2] ), .B(n18), .CI(n32), .CO(\CARRYB[2><2] ), .S(
        \SUMB[2><2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2><3] ), .B(n17), .CI(n31), .CO(\CARRYB[2><3] ), .S(
        \SUMB[2><3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2><4] ), .B(n16), .CI(n30), .CO(\CARRYB[2><4] ), .S(
        \SUMB[2><4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2><5] ), .B(n15), .CI(n29), .CO(\CARRYB[2><5] ), .S(
        \SUMB[2><5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2><6] ), .B(n14), .CI(n28), .CO(\CARRYB[2><6] ), .S(
        \SUMB[2><6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2><7] ), .B(n13), .CI(n27), .CO(\CARRYB[2><7] ), .S(
        \SUMB[2><7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2><8] ), .B(n12), .CI(n26), .CO(\CARRYB[2><8] ), .S(
        \SUMB[2><8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2><9] ), .B(n11), .CI(n25), .CO(\CARRYB[2><9] ), .S(
        \SUMB[2><9] ) );
  FA_X1 S2_2_10 ( .A(\ab[2><10] ), .B(n10), .CI(n24), .CO(\CARRYB[2><10] ), 
        .S(\SUMB[2><10] ) );
  FA_X1 S2_2_11 ( .A(\ab[2><11] ), .B(n9), .CI(n23), .CO(\CARRYB[2><11] ), .S(
        \SUMB[2><11] ) );
  FA_X1 S3_2_12 ( .A(\ab[2><12] ), .B(n37), .CI(\ab[1><13] ), .CO(
        \CARRYB[2><12] ), .S(\SUMB[2><12] ) );
  warp_generator_SHMEM_ADDR_SIZE14_DW01_add_1 FS_1 ( .A({1'b0, n2, n4, n5, n21, 
        n53, n48, n52, n47, n40, n46, n39, n38, n36, \SUMB[3><0] , \A1[0] }), 
        .B({n3, n7, n6, n8, n35, n50, n45, n49, n44, n51, n43, n42, n41, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, PRODUCT[13:2]}) );
  XOR2_X1 U2 ( .A(\CARRYB[3><12] ), .B(\ab[3><13] ), .Z(n2) );
  AND2_X1 U3 ( .A1(\CARRYB[3><12] ), .A2(\ab[3><13] ), .ZN(n3) );
  XOR2_X1 U4 ( .A(\CARRYB[3><11] ), .B(\SUMB[3><12] ), .Z(n4) );
  XOR2_X1 U5 ( .A(\CARRYB[3><10] ), .B(\SUMB[3><11] ), .Z(n5) );
  AND2_X1 U6 ( .A1(\CARRYB[3><10] ), .A2(\SUMB[3><11] ), .ZN(n6) );
  AND2_X1 U7 ( .A1(\CARRYB[3><11] ), .A2(\SUMB[3><12] ), .ZN(n7) );
  AND2_X1 U8 ( .A1(\CARRYB[3><9] ), .A2(\SUMB[3><10] ), .ZN(n8) );
  AND2_X1 U9 ( .A1(\ab[0><12] ), .A2(\ab[1><11] ), .ZN(n9) );
  AND2_X1 U10 ( .A1(\ab[0><11] ), .A2(\ab[1><10] ), .ZN(n10) );
  AND2_X1 U11 ( .A1(\ab[0><10] ), .A2(\ab[1><9] ), .ZN(n11) );
  AND2_X1 U12 ( .A1(\ab[0><9] ), .A2(\ab[1><8] ), .ZN(n12) );
  AND2_X1 U13 ( .A1(\ab[0><8] ), .A2(\ab[1><7] ), .ZN(n13) );
  AND2_X1 U14 ( .A1(\ab[0><7] ), .A2(\ab[1><6] ), .ZN(n14) );
  AND2_X1 U15 ( .A1(\ab[0><6] ), .A2(\ab[1><5] ), .ZN(n15) );
  AND2_X1 U16 ( .A1(\ab[0><5] ), .A2(\ab[1><4] ), .ZN(n16) );
  AND2_X1 U17 ( .A1(\ab[0><4] ), .A2(\ab[1><3] ), .ZN(n17) );
  AND2_X1 U18 ( .A1(\ab[0><3] ), .A2(\ab[1><2] ), .ZN(n18) );
  AND2_X1 U19 ( .A1(\ab[0><2] ), .A2(\ab[1><1] ), .ZN(n19) );
  AND2_X1 U20 ( .A1(\ab[0><1] ), .A2(\ab[1><0] ), .ZN(n20) );
  XOR2_X1 U21 ( .A(\CARRYB[3><9] ), .B(\SUMB[3><10] ), .Z(n21) );
  XOR2_X1 U22 ( .A(\ab[1><0] ), .B(\ab[0><1] ), .Z(PRODUCT[1]) );
  XOR2_X1 U23 ( .A(\ab[1><12] ), .B(\ab[0><13] ), .Z(n23) );
  XOR2_X1 U24 ( .A(\ab[1><11] ), .B(\ab[0><12] ), .Z(n24) );
  XOR2_X1 U25 ( .A(\ab[1><10] ), .B(\ab[0><11] ), .Z(n25) );
  XOR2_X1 U26 ( .A(\ab[1><9] ), .B(\ab[0><10] ), .Z(n26) );
  XOR2_X1 U27 ( .A(\ab[1><8] ), .B(\ab[0><9] ), .Z(n27) );
  XOR2_X1 U28 ( .A(\ab[1><7] ), .B(\ab[0><8] ), .Z(n28) );
  XOR2_X1 U29 ( .A(\ab[1><6] ), .B(\ab[0><7] ), .Z(n29) );
  XOR2_X1 U30 ( .A(\ab[1><5] ), .B(\ab[0><6] ), .Z(n30) );
  XOR2_X1 U31 ( .A(\ab[1><4] ), .B(\ab[0><5] ), .Z(n31) );
  XOR2_X1 U32 ( .A(\ab[1><3] ), .B(\ab[0><4] ), .Z(n32) );
  XOR2_X1 U33 ( .A(\ab[1><2] ), .B(\ab[0><3] ), .Z(n33) );
  XOR2_X1 U34 ( .A(\ab[1><1] ), .B(\ab[0><2] ), .Z(n34) );
  AND2_X1 U35 ( .A1(\CARRYB[3><8] ), .A2(\SUMB[3><9] ), .ZN(n35) );
  XOR2_X1 U36 ( .A(\CARRYB[3><0] ), .B(\SUMB[3><1] ), .Z(n36) );
  AND2_X1 U37 ( .A1(\ab[0><13] ), .A2(\ab[1><12] ), .ZN(n37) );
  XOR2_X1 U38 ( .A(\CARRYB[3><1] ), .B(\SUMB[3><2] ), .Z(n38) );
  XOR2_X1 U39 ( .A(\CARRYB[3><2] ), .B(\SUMB[3><3] ), .Z(n39) );
  XOR2_X1 U40 ( .A(\CARRYB[3><4] ), .B(\SUMB[3><5] ), .Z(n40) );
  AND2_X1 U41 ( .A1(\CARRYB[3><0] ), .A2(\SUMB[3><1] ), .ZN(n41) );
  AND2_X1 U42 ( .A1(\CARRYB[3><1] ), .A2(\SUMB[3><2] ), .ZN(n42) );
  AND2_X1 U43 ( .A1(\CARRYB[3><2] ), .A2(\SUMB[3><3] ), .ZN(n43) );
  AND2_X1 U44 ( .A1(\CARRYB[3><4] ), .A2(\SUMB[3><5] ), .ZN(n44) );
  AND2_X1 U45 ( .A1(\CARRYB[3><6] ), .A2(\SUMB[3><7] ), .ZN(n45) );
  XOR2_X1 U46 ( .A(\CARRYB[3><3] ), .B(\SUMB[3><4] ), .Z(n46) );
  XOR2_X1 U47 ( .A(\CARRYB[3><5] ), .B(\SUMB[3><6] ), .Z(n47) );
  XOR2_X1 U48 ( .A(\CARRYB[3><7] ), .B(\SUMB[3><8] ), .Z(n48) );
  AND2_X1 U49 ( .A1(\CARRYB[3><5] ), .A2(\SUMB[3><6] ), .ZN(n49) );
  AND2_X1 U50 ( .A1(\CARRYB[3><7] ), .A2(\SUMB[3><8] ), .ZN(n50) );
  AND2_X1 U51 ( .A1(\CARRYB[3><3] ), .A2(\SUMB[3><4] ), .ZN(n51) );
  XOR2_X1 U52 ( .A(\CARRYB[3><6] ), .B(\SUMB[3><7] ), .Z(n52) );
  XOR2_X1 U53 ( .A(\CARRYB[3><8] ), .B(\SUMB[3><9] ), .Z(n53) );
  INV_X1 U54 ( .A(A[1]), .ZN(n55) );
  INV_X1 U55 ( .A(A[3]), .ZN(n57) );
  INV_X1 U56 ( .A(A[0]), .ZN(n54) );
  INV_X1 U57 ( .A(A[2]), .ZN(n56) );
  INV_X1 U58 ( .A(B[1]), .ZN(n70) );
  INV_X1 U59 ( .A(B[0]), .ZN(n71) );
  INV_X1 U60 ( .A(B[2]), .ZN(n69) );
  INV_X1 U61 ( .A(B[3]), .ZN(n68) );
  INV_X1 U62 ( .A(B[6]), .ZN(n65) );
  INV_X1 U63 ( .A(B[4]), .ZN(n67) );
  INV_X1 U64 ( .A(B[5]), .ZN(n66) );
  INV_X1 U65 ( .A(B[8]), .ZN(n63) );
  INV_X1 U66 ( .A(B[7]), .ZN(n64) );
  INV_X1 U67 ( .A(B[10]), .ZN(n61) );
  INV_X1 U68 ( .A(B[9]), .ZN(n62) );
  INV_X1 U69 ( .A(B[11]), .ZN(n60) );
  INV_X1 U70 ( .A(B[12]), .ZN(n59) );
  INV_X1 U71 ( .A(B[13]), .ZN(n58) );
  NOR2_X1 U73 ( .A1(n57), .A2(n62), .ZN(\ab[3><9] ) );
  NOR2_X1 U74 ( .A1(n57), .A2(n63), .ZN(\ab[3><8] ) );
  NOR2_X1 U75 ( .A1(n57), .A2(n64), .ZN(\ab[3><7] ) );
  NOR2_X1 U76 ( .A1(n57), .A2(n65), .ZN(\ab[3><6] ) );
  NOR2_X1 U77 ( .A1(n57), .A2(n66), .ZN(\ab[3><5] ) );
  NOR2_X1 U78 ( .A1(n57), .A2(n67), .ZN(\ab[3><4] ) );
  NOR2_X1 U79 ( .A1(n57), .A2(n68), .ZN(\ab[3><3] ) );
  NOR2_X1 U80 ( .A1(n57), .A2(n69), .ZN(\ab[3><2] ) );
  NOR2_X1 U81 ( .A1(n57), .A2(n70), .ZN(\ab[3><1] ) );
  NOR2_X1 U82 ( .A1(n57), .A2(n58), .ZN(\ab[3><13] ) );
  NOR2_X1 U83 ( .A1(n57), .A2(n59), .ZN(\ab[3><12] ) );
  NOR2_X1 U84 ( .A1(n57), .A2(n60), .ZN(\ab[3><11] ) );
  NOR2_X1 U85 ( .A1(n57), .A2(n61), .ZN(\ab[3><10] ) );
  NOR2_X1 U86 ( .A1(n57), .A2(n71), .ZN(\ab[3><0] ) );
  NOR2_X1 U87 ( .A1(n62), .A2(n56), .ZN(\ab[2><9] ) );
  NOR2_X1 U88 ( .A1(n63), .A2(n56), .ZN(\ab[2><8] ) );
  NOR2_X1 U89 ( .A1(n64), .A2(n56), .ZN(\ab[2><7] ) );
  NOR2_X1 U90 ( .A1(n65), .A2(n56), .ZN(\ab[2><6] ) );
  NOR2_X1 U91 ( .A1(n66), .A2(n56), .ZN(\ab[2><5] ) );
  NOR2_X1 U92 ( .A1(n67), .A2(n56), .ZN(\ab[2><4] ) );
  NOR2_X1 U93 ( .A1(n68), .A2(n56), .ZN(\ab[2><3] ) );
  NOR2_X1 U94 ( .A1(n69), .A2(n56), .ZN(\ab[2><2] ) );
  NOR2_X1 U95 ( .A1(n70), .A2(n56), .ZN(\ab[2><1] ) );
  NOR2_X1 U96 ( .A1(n58), .A2(n56), .ZN(\ab[2><13] ) );
  NOR2_X1 U97 ( .A1(n59), .A2(n56), .ZN(\ab[2><12] ) );
  NOR2_X1 U98 ( .A1(n60), .A2(n56), .ZN(\ab[2><11] ) );
  NOR2_X1 U99 ( .A1(n61), .A2(n56), .ZN(\ab[2><10] ) );
  NOR2_X1 U100 ( .A1(n71), .A2(n56), .ZN(\ab[2><0] ) );
  NOR2_X1 U101 ( .A1(n62), .A2(n55), .ZN(\ab[1><9] ) );
  NOR2_X1 U102 ( .A1(n63), .A2(n55), .ZN(\ab[1><8] ) );
  NOR2_X1 U103 ( .A1(n64), .A2(n55), .ZN(\ab[1><7] ) );
  NOR2_X1 U104 ( .A1(n65), .A2(n55), .ZN(\ab[1><6] ) );
  NOR2_X1 U105 ( .A1(n66), .A2(n55), .ZN(\ab[1><5] ) );
  NOR2_X1 U106 ( .A1(n67), .A2(n55), .ZN(\ab[1><4] ) );
  NOR2_X1 U107 ( .A1(n68), .A2(n55), .ZN(\ab[1><3] ) );
  NOR2_X1 U108 ( .A1(n69), .A2(n55), .ZN(\ab[1><2] ) );
  NOR2_X1 U109 ( .A1(n70), .A2(n55), .ZN(\ab[1><1] ) );
  NOR2_X1 U110 ( .A1(n58), .A2(n55), .ZN(\ab[1><13] ) );
  NOR2_X1 U111 ( .A1(n59), .A2(n55), .ZN(\ab[1><12] ) );
  NOR2_X1 U112 ( .A1(n60), .A2(n55), .ZN(\ab[1><11] ) );
  NOR2_X1 U113 ( .A1(n61), .A2(n55), .ZN(\ab[1><10] ) );
  NOR2_X1 U114 ( .A1(n71), .A2(n55), .ZN(\ab[1><0] ) );
  NOR2_X1 U115 ( .A1(n62), .A2(n54), .ZN(\ab[0><9] ) );
  NOR2_X1 U116 ( .A1(n63), .A2(n54), .ZN(\ab[0><8] ) );
  NOR2_X1 U117 ( .A1(n64), .A2(n54), .ZN(\ab[0><7] ) );
  NOR2_X1 U118 ( .A1(n65), .A2(n54), .ZN(\ab[0><6] ) );
  NOR2_X1 U119 ( .A1(n66), .A2(n54), .ZN(\ab[0><5] ) );
  NOR2_X1 U120 ( .A1(n67), .A2(n54), .ZN(\ab[0><4] ) );
  NOR2_X1 U121 ( .A1(n68), .A2(n54), .ZN(\ab[0><3] ) );
  NOR2_X1 U122 ( .A1(n69), .A2(n54), .ZN(\ab[0><2] ) );
  NOR2_X1 U123 ( .A1(n70), .A2(n54), .ZN(\ab[0><1] ) );
  NOR2_X1 U124 ( .A1(n58), .A2(n54), .ZN(\ab[0><13] ) );
  NOR2_X1 U125 ( .A1(n59), .A2(n54), .ZN(\ab[0><12] ) );
  NOR2_X1 U126 ( .A1(n60), .A2(n54), .ZN(\ab[0><11] ) );
  NOR2_X1 U127 ( .A1(n61), .A2(n54), .ZN(\ab[0><10] ) );
  NOR2_X1 U128 ( .A1(n71), .A2(n54), .ZN(PRODUCT[0]) );
endmodule



module warp_generator_SHMEM_ADDR_SIZE14_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [13:1] carry;

  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .S(SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule



module warp_generator ( clk_in, host_reset, en, 
        num_blocks_in, warps_per_block_in, shmem_base_addr_in, shmem_size_in, 
        gprs_size_in, warp_pool_addr_out, warp_pool_wr_en_out, 
        warp_pool_wr_data_out, warp_state_addr_out, warp_state_wr_en_out, 
        warp_state_wr_data_out, .fence_regs_cta_id_out({
        \fence_regs_cta_id_out[31><3] , \fence_regs_cta_id_out[31><2] , 
        \fence_regs_cta_id_out[31><1] , \fence_regs_cta_id_out[31><0] , 
        \fence_regs_cta_id_out[30><3] , \fence_regs_cta_id_out[30><2] , 
        \fence_regs_cta_id_out[30><1] , \fence_regs_cta_id_out[30><0] , 
        \fence_regs_cta_id_out[29><3] , \fence_regs_cta_id_out[29><2] , 
        \fence_regs_cta_id_out[29><1] , \fence_regs_cta_id_out[29><0] , 
        \fence_regs_cta_id_out[28><3] , \fence_regs_cta_id_out[28><2] , 
        \fence_regs_cta_id_out[28><1] , \fence_regs_cta_id_out[28><0] , 
        \fence_regs_cta_id_out[27><3] , \fence_regs_cta_id_out[27><2] , 
        \fence_regs_cta_id_out[27><1] , \fence_regs_cta_id_out[27><0] , 
        \fence_regs_cta_id_out[26><3] , \fence_regs_cta_id_out[26><2] , 
        \fence_regs_cta_id_out[26><1] , \fence_regs_cta_id_out[26><0] , 
        \fence_regs_cta_id_out[25><3] , \fence_regs_cta_id_out[25><2] , 
        \fence_regs_cta_id_out[25><1] , \fence_regs_cta_id_out[25><0] , 
        \fence_regs_cta_id_out[24><3] , \fence_regs_cta_id_out[24><2] , 
        \fence_regs_cta_id_out[24><1] , \fence_regs_cta_id_out[24><0] , 
        \fence_regs_cta_id_out[23><3] , \fence_regs_cta_id_out[23><2] , 
        \fence_regs_cta_id_out[23><1] , \fence_regs_cta_id_out[23><0] , 
        \fence_regs_cta_id_out[22><3] , \fence_regs_cta_id_out[22><2] , 
        \fence_regs_cta_id_out[22><1] , \fence_regs_cta_id_out[22><0] , 
        \fence_regs_cta_id_out[21><3] , \fence_regs_cta_id_out[21><2] , 
        \fence_regs_cta_id_out[21><1] , \fence_regs_cta_id_out[21><0] , 
        \fence_regs_cta_id_out[20><3] , \fence_regs_cta_id_out[20><2] , 
        \fence_regs_cta_id_out[20><1] , \fence_regs_cta_id_out[20><0] , 
        \fence_regs_cta_id_out[19><3] , \fence_regs_cta_id_out[19><2] , 
        \fence_regs_cta_id_out[19><1] , \fence_regs_cta_id_out[19><0] , 
        \fence_regs_cta_id_out[18><3] , \fence_regs_cta_id_out[18><2] , 
        \fence_regs_cta_id_out[18><1] , \fence_regs_cta_id_out[18><0] , 
        \fence_regs_cta_id_out[17><3] , \fence_regs_cta_id_out[17><2] , 
        \fence_regs_cta_id_out[17><1] , \fence_regs_cta_id_out[17><0] , 
        \fence_regs_cta_id_out[16><3] , \fence_regs_cta_id_out[16><2] , 
        \fence_regs_cta_id_out[16><1] , \fence_regs_cta_id_out[16><0] , 
        \fence_regs_cta_id_out[15><3] , \fence_regs_cta_id_out[15><2] , 
        \fence_regs_cta_id_out[15><1] , \fence_regs_cta_id_out[15><0] , 
        \fence_regs_cta_id_out[14><3] , \fence_regs_cta_id_out[14><2] , 
        \fence_regs_cta_id_out[14><1] , \fence_regs_cta_id_out[14><0] , 
        \fence_regs_cta_id_out[13><3] , \fence_regs_cta_id_out[13><2] , 
        \fence_regs_cta_id_out[13><1] , \fence_regs_cta_id_out[13><0] , 
        \fence_regs_cta_id_out[12><3] , \fence_regs_cta_id_out[12><2] , 
        \fence_regs_cta_id_out[12><1] , \fence_regs_cta_id_out[12><0] , 
        \fence_regs_cta_id_out[11><3] , \fence_regs_cta_id_out[11><2] , 
        \fence_regs_cta_id_out[11><1] , \fence_regs_cta_id_out[11><0] , 
        \fence_regs_cta_id_out[10><3] , \fence_regs_cta_id_out[10><2] , 
        \fence_regs_cta_id_out[10><1] , \fence_regs_cta_id_out[10><0] , 
        \fence_regs_cta_id_out[9><3] , \fence_regs_cta_id_out[9><2] , 
        \fence_regs_cta_id_out[9><1] , \fence_regs_cta_id_out[9><0] , 
        \fence_regs_cta_id_out[8><3] , \fence_regs_cta_id_out[8><2] , 
        \fence_regs_cta_id_out[8><1] , \fence_regs_cta_id_out[8><0] , 
        \fence_regs_cta_id_out[7><3] , \fence_regs_cta_id_out[7><2] , 
        \fence_regs_cta_id_out[7><1] , \fence_regs_cta_id_out[7><0] , 
        \fence_regs_cta_id_out[6><3] , \fence_regs_cta_id_out[6><2] , 
        \fence_regs_cta_id_out[6><1] , \fence_regs_cta_id_out[6><0] , 
        \fence_regs_cta_id_out[5><3] , \fence_regs_cta_id_out[5><2] , 
        \fence_regs_cta_id_out[5><1] , \fence_regs_cta_id_out[5><0] , 
        \fence_regs_cta_id_out[4><3] , \fence_regs_cta_id_out[4><2] , 
        \fence_regs_cta_id_out[4><1] , \fence_regs_cta_id_out[4><0] , 
        \fence_regs_cta_id_out[3><3] , \fence_regs_cta_id_out[3><2] , 
        \fence_regs_cta_id_out[3><1] , \fence_regs_cta_id_out[3><0] , 
        \fence_regs_cta_id_out[2><3] , \fence_regs_cta_id_out[2><2] , 
        \fence_regs_cta_id_out[2><1] , \fence_regs_cta_id_out[2><0] , 
        \fence_regs_cta_id_out[1><3] , \fence_regs_cta_id_out[1><2] , 
        \fence_regs_cta_id_out[1><1] , \fence_regs_cta_id_out[1><0] , 
        \fence_regs_cta_id_out[0><3] , \fence_regs_cta_id_out[0><2] , 
        \fence_regs_cta_id_out[0><1] , \fence_regs_cta_id_out[0><0] }), 
        fence_regs_cta_id_ld, fence_regs_fence_en_out, fence_regs_fence_en_ld, 
        num_warps_out, warp_gen_done );
  input [3:0] num_blocks_in;
  input [5:0] warps_per_block_in;
  input [31:0] shmem_base_addr_in;
  input [31:0] shmem_size_in;
  input [8:0] gprs_size_in;
  output [4:0] warp_pool_addr_out;
  output [127:0] warp_pool_wr_data_out;
  output [4:0] warp_state_addr_out;
  output [1:0] warp_state_wr_data_out;
  output [31:0] fence_regs_cta_id_ld;
  output [31:0] fence_regs_fence_en_out;
  output [31:0] fence_regs_fence_en_ld;
  output [4:0] num_warps_out;
  input clk_in, host_reset, en;
  output warp_pool_wr_en_out, warp_state_wr_en_out,
         \fence_regs_cta_id_out[31><3] , \fence_regs_cta_id_out[31><2] ,
         \fence_regs_cta_id_out[31><1] , \fence_regs_cta_id_out[31><0] ,
         \fence_regs_cta_id_out[30><3] , \fence_regs_cta_id_out[30><2] ,
         \fence_regs_cta_id_out[30><1] , \fence_regs_cta_id_out[30><0] ,
         \fence_regs_cta_id_out[29><3] , \fence_regs_cta_id_out[29><2] ,
         \fence_regs_cta_id_out[29><1] , \fence_regs_cta_id_out[29><0] ,
         \fence_regs_cta_id_out[28><3] , \fence_regs_cta_id_out[28><2] ,
         \fence_regs_cta_id_out[28><1] , \fence_regs_cta_id_out[28><0] ,
         \fence_regs_cta_id_out[27><3] , \fence_regs_cta_id_out[27><2] ,
         \fence_regs_cta_id_out[27><1] , \fence_regs_cta_id_out[27><0] ,
         \fence_regs_cta_id_out[26><3] , \fence_regs_cta_id_out[26><2] ,
         \fence_regs_cta_id_out[26><1] , \fence_regs_cta_id_out[26><0] ,
         \fence_regs_cta_id_out[25><3] , \fence_regs_cta_id_out[25><2] ,
         \fence_regs_cta_id_out[25><1] , \fence_regs_cta_id_out[25><0] ,
         \fence_regs_cta_id_out[24><3] , \fence_regs_cta_id_out[24><2] ,
         \fence_regs_cta_id_out[24><1] , \fence_regs_cta_id_out[24><0] ,
         \fence_regs_cta_id_out[23><3] , \fence_regs_cta_id_out[23><2] ,
         \fence_regs_cta_id_out[23><1] , \fence_regs_cta_id_out[23><0] ,
         \fence_regs_cta_id_out[22><3] , \fence_regs_cta_id_out[22><2] ,
         \fence_regs_cta_id_out[22><1] , \fence_regs_cta_id_out[22><0] ,
         \fence_regs_cta_id_out[21><3] , \fence_regs_cta_id_out[21><2] ,
         \fence_regs_cta_id_out[21><1] , \fence_regs_cta_id_out[21><0] ,
         \fence_regs_cta_id_out[20><3] , \fence_regs_cta_id_out[20><2] ,
         \fence_regs_cta_id_out[20><1] , \fence_regs_cta_id_out[20><0] ,
         \fence_regs_cta_id_out[19><3] , \fence_regs_cta_id_out[19><2] ,
         \fence_regs_cta_id_out[19><1] , \fence_regs_cta_id_out[19><0] ,
         \fence_regs_cta_id_out[18><3] , \fence_regs_cta_id_out[18><2] ,
         \fence_regs_cta_id_out[18><1] , \fence_regs_cta_id_out[18><0] ,
         \fence_regs_cta_id_out[17><3] , \fence_regs_cta_id_out[17><2] ,
         \fence_regs_cta_id_out[17><1] , \fence_regs_cta_id_out[17><0] ,
         \fence_regs_cta_id_out[16><3] , \fence_regs_cta_id_out[16><2] ,
         \fence_regs_cta_id_out[16><1] , \fence_regs_cta_id_out[16><0] ,
         \fence_regs_cta_id_out[15><3] , \fence_regs_cta_id_out[15><2] ,
         \fence_regs_cta_id_out[15><1] , \fence_regs_cta_id_out[15><0] ,
         \fence_regs_cta_id_out[14><3] , \fence_regs_cta_id_out[14><2] ,
         \fence_regs_cta_id_out[14><1] , \fence_regs_cta_id_out[14><0] ,
         \fence_regs_cta_id_out[13><3] , \fence_regs_cta_id_out[13><2] ,
         \fence_regs_cta_id_out[13><1] , \fence_regs_cta_id_out[13><0] ,
         \fence_regs_cta_id_out[12><3] , \fence_regs_cta_id_out[12><2] ,
         \fence_regs_cta_id_out[12><1] , \fence_regs_cta_id_out[12><0] ,
         \fence_regs_cta_id_out[11><3] , \fence_regs_cta_id_out[11><2] ,
         \fence_regs_cta_id_out[11><1] , \fence_regs_cta_id_out[11><0] ,
         \fence_regs_cta_id_out[10><3] , \fence_regs_cta_id_out[10><2] ,
         \fence_regs_cta_id_out[10><1] , \fence_regs_cta_id_out[10><0] ,
         \fence_regs_cta_id_out[9><3] , \fence_regs_cta_id_out[9><2] ,
         \fence_regs_cta_id_out[9><1] , \fence_regs_cta_id_out[9><0] ,
         \fence_regs_cta_id_out[8><3] , \fence_regs_cta_id_out[8><2] ,
         \fence_regs_cta_id_out[8><1] , \fence_regs_cta_id_out[8><0] ,
         \fence_regs_cta_id_out[7><3] , \fence_regs_cta_id_out[7><2] ,
         \fence_regs_cta_id_out[7><1] , \fence_regs_cta_id_out[7><0] ,
         \fence_regs_cta_id_out[6><3] , \fence_regs_cta_id_out[6><2] ,
         \fence_regs_cta_id_out[6><1] , \fence_regs_cta_id_out[6><0] ,
         \fence_regs_cta_id_out[5><3] , \fence_regs_cta_id_out[5><2] ,
         \fence_regs_cta_id_out[5><1] , \fence_regs_cta_id_out[5><0] ,
         \fence_regs_cta_id_out[4><3] , \fence_regs_cta_id_out[4><2] ,
         \fence_regs_cta_id_out[4><1] , \fence_regs_cta_id_out[4><0] ,
         \fence_regs_cta_id_out[3><3] , \fence_regs_cta_id_out[3><2] ,
         \fence_regs_cta_id_out[3><1] , \fence_regs_cta_id_out[3><0] ,
         \fence_regs_cta_id_out[2><3] , \fence_regs_cta_id_out[2><2] ,
         \fence_regs_cta_id_out[2><1] , \fence_regs_cta_id_out[2><0] ,
         \fence_regs_cta_id_out[1><3] , \fence_regs_cta_id_out[1><2] ,
         \fence_regs_cta_id_out[1><1] , \fence_regs_cta_id_out[1><0] ,
         \fence_regs_cta_id_out[0><3] , \fence_regs_cta_id_out[0><2] ,
         \fence_regs_cta_id_out[0><1] , \fence_regs_cta_id_out[0><0] ,
         warp_gen_done;
  wire   warp_id_calc_en_i, N62, N78, N79, N80, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N254, N255, N256, N257, N863, N864, N865, N866,
         N867, N868, N869, N870, N871, N872, N873, N874, N875, N876, N877,
         N878, N879, N880, N881, N882, N883, N884, N885, N886, N887, N888,
         N889, N890, N891, N892, N893, N894, n40, n41, n42, n43, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n141, n142, n143, n145,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67,
         N66, N65, N64, \add_155/carry[4] , \add_155/carry[3] ,
         \add_155/carry[2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n144, n146, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n272, n273,
         n274, n275, n276, n277, n278, n279, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876;
  wire   [3:0] block_num_cnt;
  wire   [11:0] warps_per_block_cnt;
  wire   [3:0] block_num_i;
  wire   [4:0] warp_num_i;
  wire   [2:0] warp_generator_state_machine;
  wire   [13:0] shmem_addr_i;
  wire   [4:0] warp_id_o;
  wire   [4:0] warp_id_addr;
  wire   [8:0] gprs_base_addr_o;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign warp_pool_wr_data_out[127] = 1'b0;
  assign warp_pool_wr_data_out[126] = 1'b0;
  assign warp_pool_wr_data_out[125] = 1'b0;
  assign warp_pool_wr_data_out[124] = 1'b0;
  assign warp_pool_wr_data_out[96] = 1'b0;
  assign warp_pool_wr_data_out[95] = 1'b0;
  assign warp_pool_wr_data_out[94] = 1'b0;
  assign warp_pool_wr_data_out[93] = 1'b0;
  assign warp_pool_wr_data_out[92] = 1'b0;
  assign warp_pool_wr_data_out[91] = 1'b0;
  assign warp_pool_wr_data_out[90] = 1'b0;
  assign warp_pool_wr_data_out[89] = 1'b0;
  assign warp_pool_wr_data_out[88] = 1'b0;
  assign warp_pool_wr_data_out[87] = 1'b0;
  assign warp_pool_wr_data_out[86] = 1'b0;
  assign warp_pool_wr_data_out[85] = 1'b0;
  assign warp_pool_wr_data_out[84] = 1'b0;
  assign warp_pool_wr_data_out[83] = 1'b0;
  assign warp_pool_wr_data_out[82] = 1'b0;
  assign warp_pool_wr_data_out[81] = 1'b0;
  assign warp_pool_wr_data_out[80] = 1'b0;
  assign warp_pool_wr_data_out[79] = 1'b0;
  assign warp_pool_wr_data_out[78] = 1'b0;
  assign warp_pool_wr_data_out[77] = 1'b0;
  assign warp_pool_wr_data_out[76] = 1'b0;
  assign warp_pool_wr_data_out[75] = 1'b0;
  assign warp_pool_wr_data_out[74] = 1'b0;
  assign warp_pool_wr_data_out[73] = 1'b0;
  assign warp_pool_wr_data_out[72] = 1'b0;
  assign warp_pool_wr_data_out[71] = 1'b0;
  assign warp_pool_wr_data_out[70] = 1'b0;
  assign warp_pool_wr_data_out[69] = 1'b0;
  assign warp_pool_wr_data_out[68] = 1'b0;
  assign warp_pool_wr_data_out[67] = 1'b0;
  assign warp_pool_wr_data_out[66] = 1'b0;
  assign warp_pool_wr_data_out[65] = 1'b0;
  assign warp_pool_wr_data_out[64] = 1'b0;
  assign warp_state_wr_data_out[1] = 1'b0;
  assign warp_state_wr_data_out[0] = 1'b0;
  assign fence_regs_fence_en_out[31] = 1'b0;
  assign fence_regs_fence_en_out[30] = 1'b0;
  assign fence_regs_fence_en_out[29] = 1'b0;
  assign fence_regs_fence_en_out[28] = 1'b0;
  assign fence_regs_fence_en_out[27] = 1'b0;
  assign fence_regs_fence_en_out[26] = 1'b0;
  assign fence_regs_fence_en_out[25] = 1'b0;
  assign fence_regs_fence_en_out[24] = 1'b0;
  assign fence_regs_fence_en_out[23] = 1'b0;
  assign fence_regs_fence_en_out[22] = 1'b0;
  assign fence_regs_fence_en_out[21] = 1'b0;
  assign fence_regs_fence_en_out[20] = 1'b0;
  assign fence_regs_fence_en_out[19] = 1'b0;
  assign fence_regs_fence_en_out[18] = 1'b0;
  assign fence_regs_fence_en_out[17] = 1'b0;
  assign fence_regs_fence_en_out[16] = 1'b0;
  assign fence_regs_fence_en_out[15] = 1'b0;
  assign fence_regs_fence_en_out[14] = 1'b0;
  assign fence_regs_fence_en_out[13] = 1'b0;
  assign fence_regs_fence_en_out[12] = 1'b0;
  assign fence_regs_fence_en_out[11] = 1'b0;
  assign fence_regs_fence_en_out[10] = 1'b0;
  assign fence_regs_fence_en_out[9] = 1'b0;
  assign fence_regs_fence_en_out[8] = 1'b0;
  assign fence_regs_fence_en_out[7] = 1'b0;
  assign fence_regs_fence_en_out[6] = 1'b0;
  assign fence_regs_fence_en_out[5] = 1'b0;
  assign fence_regs_fence_en_out[4] = 1'b0;
  assign fence_regs_fence_en_out[3] = 1'b0;
  assign fence_regs_fence_en_out[2] = 1'b0;
  assign fence_regs_fence_en_out[1] = 1'b0;
  assign fence_regs_fence_en_out[0] = 1'b0;

  DFFR_X1 \warp_generator_state_machine_reg[0]  ( .D(n815), .CK(clk_in), .RN(
        n121), .Q(warp_generator_state_machine[0]), .QN(n202) );
  DFFR_X1 \warp_generator_state_machine_reg[1]  ( .D(n814), .CK(clk_in), .RN(
        n121), .Q(warp_generator_state_machine[1]), .QN(n201) );
  DFFR_X1 \warps_per_block_cnt_reg[11]  ( .D(n277), .CK(clk_in), .RN(n121), 
        .Q(warps_per_block_cnt[11]) );
  DFFR_X1 \warps_per_block_cnt_reg[0]  ( .D(n278), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[0]), .QN(n151) );
  DFFR_X1 \warps_per_block_cnt_reg[1]  ( .D(n279), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[1]), .QN(n150) );
  DFFR_X1 \warps_per_block_cnt_reg[2]  ( .D(n816), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[2]), .QN(n149) );
  DFFR_X1 \warps_per_block_cnt_reg[3]  ( .D(n817), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[3]), .QN(n148) );
  DFFR_X1 \warps_per_block_cnt_reg[4]  ( .D(n818), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[4]), .QN(n147) );
  DFFR_X1 \warps_per_block_cnt_reg[5]  ( .D(n819), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[5]), .QN(n2) );
  DFFR_X1 \warps_per_block_cnt_reg[6]  ( .D(n820), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[6]) );
  DFFR_X1 \warps_per_block_cnt_reg[7]  ( .D(n821), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[7]) );
  DFFR_X1 \warps_per_block_cnt_reg[8]  ( .D(n822), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[8]) );
  DFFR_X1 \warps_per_block_cnt_reg[9]  ( .D(n823), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[9]) );
  DFFR_X1 \warps_per_block_cnt_reg[10]  ( .D(n824), .CK(clk_in), .RN(n121), 
        .Q(warps_per_block_cnt[10]) );
  DFFR_X1 \block_num_cnt_reg[0]  ( .D(n810), .CK(clk_in), .RN(n121), .Q(
        block_num_cnt[0]), .QN(n145) );
  DFFR_X1 \block_num_cnt_reg[1]  ( .D(n811), .CK(clk_in), .RN(n121), .Q(
        block_num_cnt[1]), .QN(n143) );
  DFFR_X1 \block_num_cnt_reg[2]  ( .D(n809), .CK(clk_in), .RN(n121), .Q(
        block_num_cnt[2]), .QN(n142) );
  DFFR_X1 \block_num_cnt_reg[3]  ( .D(n808), .CK(clk_in), .RN(n121), .Q(
        block_num_cnt[3]), .QN(n141) );
  DFFR_X1 \warp_generator_state_machine_reg[2]  ( .D(n197), .CK(clk_in), .RN(
        n122), .Q(warp_generator_state_machine[2]), .QN(n200) );
  DFFR_X1 warp_state_wr_en_out_reg ( .D(n812), .CK(clk_in), .RN(n122), .Q(
        warp_state_wr_en_out) );
  DFFR_X1 warp_pool_wr_en_out_reg ( .D(n813), .CK(clk_in), .RN(n122), .Q(
        warp_pool_wr_en_out) );
  DFFR_X1 \warp_pool_wr_data_out_reg[0]  ( .D(n733), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[0]), .QN(n116) );
  DFFR_X1 \warp_pool_wr_data_out_reg[63]  ( .D(n734), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[63]), .QN(n53) );
  DFFR_X1 \warp_pool_wr_data_out_reg[62]  ( .D(n735), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[62]), .QN(n54) );
  DFFR_X1 \warp_pool_wr_data_out_reg[61]  ( .D(n736), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[61]), .QN(n55) );
  DFFR_X1 \warp_pool_wr_data_out_reg[60]  ( .D(n737), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[60]), .QN(n56) );
  DFFR_X1 \warp_pool_wr_data_out_reg[59]  ( .D(n738), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[59]), .QN(n57) );
  DFFR_X1 \warp_pool_wr_data_out_reg[58]  ( .D(n739), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[58]), .QN(n58) );
  DFFR_X1 \warp_pool_wr_data_out_reg[57]  ( .D(n740), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[57]), .QN(n59) );
  DFFR_X1 \warp_pool_wr_data_out_reg[56]  ( .D(n741), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[56]), .QN(n60) );
  DFFR_X1 \warp_pool_wr_data_out_reg[55]  ( .D(n742), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[55]), .QN(n61) );
  DFFR_X1 \warp_pool_wr_data_out_reg[54]  ( .D(n743), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[54]), .QN(n62) );
  DFFR_X1 \warp_pool_wr_data_out_reg[53]  ( .D(n744), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[53]), .QN(n63) );
  DFFR_X1 \warp_pool_wr_data_out_reg[52]  ( .D(n745), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[52]), .QN(n64) );
  DFFR_X1 \warp_pool_wr_data_out_reg[51]  ( .D(n746), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[51]), .QN(n65) );
  DFFR_X1 \warp_pool_wr_data_out_reg[50]  ( .D(n747), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[50]), .QN(n66) );
  DFFR_X1 \warp_pool_wr_data_out_reg[49]  ( .D(n748), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[49]), .QN(n67) );
  DFFR_X1 \warp_pool_wr_data_out_reg[48]  ( .D(n749), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[48]), .QN(n68) );
  DFFR_X1 \warp_pool_wr_data_out_reg[47]  ( .D(n750), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[47]), .QN(n69) );
  DFFR_X1 \warp_pool_wr_data_out_reg[46]  ( .D(n751), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[46]), .QN(n70) );
  DFFR_X1 \warp_pool_wr_data_out_reg[45]  ( .D(n752), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[45]), .QN(n71) );
  DFFR_X1 \warp_pool_wr_data_out_reg[44]  ( .D(n753), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[44]), .QN(n72) );
  DFFR_X1 \warp_pool_wr_data_out_reg[43]  ( .D(n754), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[43]), .QN(n73) );
  DFFR_X1 \warp_pool_wr_data_out_reg[42]  ( .D(n755), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[42]), .QN(n74) );
  DFFR_X1 \warp_pool_wr_data_out_reg[41]  ( .D(n756), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[41]), .QN(n75) );
  DFFR_X1 \warp_pool_wr_data_out_reg[40]  ( .D(n757), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[40]), .QN(n76) );
  DFFR_X1 \warp_pool_wr_data_out_reg[39]  ( .D(n758), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[39]), .QN(n77) );
  DFFR_X1 \warp_pool_wr_data_out_reg[38]  ( .D(n759), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[38]), .QN(n78) );
  DFFR_X1 \warp_pool_wr_data_out_reg[37]  ( .D(n760), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[37]), .QN(n79) );
  DFFR_X1 \warp_pool_wr_data_out_reg[36]  ( .D(n761), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[36]), .QN(n80) );
  DFFR_X1 \warp_pool_wr_data_out_reg[35]  ( .D(n762), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[35]), .QN(n81) );
  DFFR_X1 \warp_pool_wr_data_out_reg[34]  ( .D(n763), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[34]), .QN(n82) );
  DFFR_X1 \warp_pool_wr_data_out_reg[33]  ( .D(n764), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[33]), .QN(n83) );
  DFFR_X1 \warp_pool_wr_data_out_reg[32]  ( .D(n765), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[32]), .QN(n84) );
  DFFR_X1 \warp_pool_wr_data_out_reg[31]  ( .D(n766), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[31]), .QN(n85) );
  DFFR_X1 \warp_pool_wr_data_out_reg[30]  ( .D(n767), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[30]), .QN(n86) );
  DFFR_X1 \warp_pool_wr_data_out_reg[29]  ( .D(n768), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[29]), .QN(n87) );
  DFFR_X1 \warp_pool_wr_data_out_reg[28]  ( .D(n769), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[28]), .QN(n88) );
  DFFR_X1 \warp_pool_wr_data_out_reg[27]  ( .D(n770), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[27]), .QN(n89) );
  DFFR_X1 \warp_pool_wr_data_out_reg[26]  ( .D(n771), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[26]), .QN(n90) );
  DFFR_X1 \warp_pool_wr_data_out_reg[25]  ( .D(n772), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[25]), .QN(n91) );
  DFFR_X1 \warp_pool_wr_data_out_reg[24]  ( .D(n773), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[24]), .QN(n92) );
  DFFR_X1 \warp_pool_wr_data_out_reg[23]  ( .D(n774), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[23]), .QN(n93) );
  DFFR_X1 \warp_pool_wr_data_out_reg[22]  ( .D(n775), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[22]), .QN(n94) );
  DFFR_X1 \warp_pool_wr_data_out_reg[21]  ( .D(n776), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[21]), .QN(n95) );
  DFFR_X1 \warp_pool_wr_data_out_reg[20]  ( .D(n777), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[20]), .QN(n96) );
  DFFR_X1 \warp_pool_wr_data_out_reg[19]  ( .D(n778), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[19]), .QN(n97) );
  DFFR_X1 \warp_pool_wr_data_out_reg[18]  ( .D(n779), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[18]), .QN(n98) );
  DFFR_X1 \warp_pool_wr_data_out_reg[17]  ( .D(n780), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[17]), .QN(n99) );
  DFFR_X1 \warp_pool_wr_data_out_reg[16]  ( .D(n781), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[16]), .QN(n100) );
  DFFR_X1 \warp_pool_wr_data_out_reg[15]  ( .D(n782), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[15]), .QN(n101) );
  DFFR_X1 \warp_pool_wr_data_out_reg[14]  ( .D(n783), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[14]), .QN(n102) );
  DFFR_X1 \warp_pool_wr_data_out_reg[13]  ( .D(n784), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[13]), .QN(n103) );
  DFFR_X1 \warp_pool_wr_data_out_reg[12]  ( .D(n785), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[12]), .QN(n104) );
  DFFR_X1 \warp_pool_wr_data_out_reg[11]  ( .D(n786), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[11]), .QN(n105) );
  DFFR_X1 \warp_pool_wr_data_out_reg[10]  ( .D(n787), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[10]), .QN(n106) );
  DFFR_X1 \warp_pool_wr_data_out_reg[9]  ( .D(n788), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[9]), .QN(n107) );
  DFFR_X1 \warp_pool_wr_data_out_reg[8]  ( .D(n789), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[8]), .QN(n108) );
  DFFR_X1 \warp_pool_wr_data_out_reg[7]  ( .D(n790), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[7]), .QN(n109) );
  DFFR_X1 \warp_pool_wr_data_out_reg[6]  ( .D(n791), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[6]), .QN(n110) );
  DFFR_X1 \warp_pool_wr_data_out_reg[5]  ( .D(n792), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[5]), .QN(n111) );
  DFFR_X1 \warp_pool_wr_data_out_reg[4]  ( .D(n793), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[4]), .QN(n112) );
  DFFR_X1 \warp_pool_wr_data_out_reg[3]  ( .D(n794), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[3]), .QN(n113) );
  DFFR_X1 \warp_pool_wr_data_out_reg[2]  ( .D(n795), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[2]), .QN(n114) );
  DFFR_X1 \warp_pool_wr_data_out_reg[1]  ( .D(n796), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[1]), .QN(n115) );
  DFFR_X1 \warp_num_i_reg[0]  ( .D(n802), .CK(clk_in), .RN(n125), .Q(
        warp_num_i[0]) );
  DFFR_X1 \warp_num_i_reg[1]  ( .D(n803), .CK(clk_in), .RN(n125), .Q(
        warp_num_i[1]) );
  DFFR_X1 \warp_num_i_reg[2]  ( .D(n804), .CK(clk_in), .RN(n125), .Q(
        warp_num_i[2]) );
  DFFR_X1 \warp_num_i_reg[3]  ( .D(n805), .CK(clk_in), .RN(n125), .Q(
        warp_num_i[3]) );
  DFFR_X1 \warp_num_i_reg[4]  ( .D(n806), .CK(clk_in), .RN(n125), .Q(
        warp_num_i[4]) );
  DFFR_X1 warp_id_calc_en_i_reg ( .D(n798), .CK(clk_in), .RN(n125), .Q(
        warp_id_calc_en_i), .QN(n156) );
  DFFR_X1 \block_num_i_reg[1]  ( .D(n799), .CK(clk_in), .RN(n125), .Q(
        block_num_i[1]), .QN(n154) );
  DFFR_X1 \warp_pool_wr_data_out_reg[107]  ( .D(n731), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[107]), .QN(n42) );
  DFFR_X1 \block_num_i_reg[2]  ( .D(n800), .CK(clk_in), .RN(n125), .Q(
        block_num_i[2]), .QN(n153) );
  DFFR_X1 \warp_pool_wr_data_out_reg[108]  ( .D(n730), .CK(clk_in), .RN(n126), 
        .Q(warp_pool_wr_data_out[108]), .QN(n41) );
  DFFR_X1 \block_num_i_reg[3]  ( .D(n801), .CK(clk_in), .RN(n126), .Q(
        block_num_i[3]), .QN(n152) );
  DFFR_X1 \warp_pool_wr_data_out_reg[109]  ( .D(n729), .CK(clk_in), .RN(n126), 
        .Q(warp_pool_wr_data_out[109]), .QN(n40) );
  DFFR_X1 \block_num_i_reg[0]  ( .D(n807), .CK(clk_in), .RN(n126), .Q(
        block_num_i[0]), .QN(n155) );
  DFFR_X1 \warp_state_addr_out_reg[0]  ( .D(n182), .CK(clk_in), .RN(n126), .Q(
        warp_state_addr_out[0]) );
  DFFR_X1 \warp_pool_addr_out_reg[0]  ( .D(n181), .CK(clk_in), .RN(n126), .Q(
        warp_pool_addr_out[0]) );
  DFFR_X1 \warp_state_addr_out_reg[1]  ( .D(n177), .CK(clk_in), .RN(n126), .Q(
        warp_state_addr_out[1]) );
  DFFR_X1 \warp_pool_addr_out_reg[1]  ( .D(n176), .CK(clk_in), .RN(n126), .Q(
        warp_pool_addr_out[1]) );
  DFFR_X1 \warp_state_addr_out_reg[2]  ( .D(n173), .CK(clk_in), .RN(n126), .Q(
        warp_state_addr_out[2]) );
  DFFR_X1 \warp_pool_addr_out_reg[2]  ( .D(n172), .CK(clk_in), .RN(n126), .Q(
        warp_pool_addr_out[2]) );
  DFFR_X1 \warp_state_addr_out_reg[3]  ( .D(n169), .CK(clk_in), .RN(n126), .Q(
        warp_state_addr_out[3]) );
  DFFR_X1 \warp_pool_addr_out_reg[3]  ( .D(n168), .CK(clk_in), .RN(n126), .Q(
        warp_pool_addr_out[3]) );
  DFFR_X1 \warp_state_addr_out_reg[4]  ( .D(n165), .CK(clk_in), .RN(n126), .Q(
        warp_state_addr_out[4]) );
  DFFR_X1 \warp_pool_addr_out_reg[4]  ( .D(n164), .CK(clk_in), .RN(n126), .Q(
        warp_pool_addr_out[4]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[97]  ( .D(n178), .CK(clk_in), .RN(n126), 
        .Q(warp_pool_wr_data_out[97]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[98]  ( .D(n161), .CK(clk_in), .RN(n126), 
        .Q(warp_pool_wr_data_out[98]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[99]  ( .D(n160), .CK(clk_in), .RN(n126), 
        .Q(warp_pool_wr_data_out[99]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[100]  ( .D(n159), .CK(clk_in), .RN(n126), 
        .Q(warp_pool_wr_data_out[100]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[101]  ( .D(n158), .CK(clk_in), .RN(n126), 
        .Q(warp_pool_wr_data_out[101]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[102]  ( .D(n157), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[102]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[103]  ( .D(n146), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[103]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[104]  ( .D(n144), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[104]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[105]  ( .D(n140), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[105]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[106]  ( .D(n732), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[106]), .QN(n43) );
  DFFR_X1 warp_gen_done_reg ( .D(n797), .CK(clk_in), .RN(n127), .Q(
        warp_gen_done) );
  DFFR_X1 \num_warps_out_reg[1]  ( .D(n174), .CK(clk_in), .RN(n127), .Q(
        num_warps_out[1]) );
  DFFR_X1 \num_warps_out_reg[2]  ( .D(n170), .CK(clk_in), .RN(n127), .Q(
        num_warps_out[2]) );
  DFFR_X1 \num_warps_out_reg[3]  ( .D(n166), .CK(clk_in), .RN(n127), .Q(
        num_warps_out[3]) );
  DFFR_X1 \num_warps_out_reg[4]  ( .D(n162), .CK(clk_in), .RN(n127), .Q(
        num_warps_out[4]) );
  DFFR_X1 \num_warps_out_reg[0]  ( .D(n179), .CK(clk_in), .RN(n127), .Q(
        num_warps_out[0]) );
  DFF_X1 \shmem_addr_i_reg[13]  ( .D(n183), .CK(clk_in), .Q(shmem_addr_i[13])
         );
  DFFR_X1 \warp_pool_wr_data_out_reg[123]  ( .D(n858), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[123]) );
  DFF_X1 \shmem_addr_i_reg[12]  ( .D(n184), .CK(clk_in), .Q(shmem_addr_i[12])
         );
  DFFR_X1 \warp_pool_wr_data_out_reg[122]  ( .D(n859), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[122]) );
  DFF_X1 \shmem_addr_i_reg[11]  ( .D(n185), .CK(clk_in), .Q(shmem_addr_i[11])
         );
  DFFR_X1 \warp_pool_wr_data_out_reg[121]  ( .D(n860), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[121]) );
  DFF_X1 \shmem_addr_i_reg[10]  ( .D(n186), .CK(clk_in), .Q(shmem_addr_i[10])
         );
  DFFR_X1 \warp_pool_wr_data_out_reg[120]  ( .D(n861), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[120]) );
  DFF_X1 \shmem_addr_i_reg[9]  ( .D(n187), .CK(clk_in), .Q(shmem_addr_i[9]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[119]  ( .D(n862), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[119]) );
  DFF_X1 \shmem_addr_i_reg[8]  ( .D(n188), .CK(clk_in), .Q(shmem_addr_i[8]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[118]  ( .D(n863), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[118]) );
  DFF_X1 \shmem_addr_i_reg[7]  ( .D(n189), .CK(clk_in), .Q(shmem_addr_i[7]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[117]  ( .D(n864), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[117]) );
  DFF_X1 \shmem_addr_i_reg[6]  ( .D(n190), .CK(clk_in), .Q(shmem_addr_i[6]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[116]  ( .D(n865), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[116]) );
  DFF_X1 \shmem_addr_i_reg[5]  ( .D(n191), .CK(clk_in), .Q(shmem_addr_i[5]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[115]  ( .D(n866), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[115]) );
  DFF_X1 \shmem_addr_i_reg[4]  ( .D(n192), .CK(clk_in), .Q(shmem_addr_i[4]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[114]  ( .D(n867), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[114]) );
  DFF_X1 \shmem_addr_i_reg[3]  ( .D(n193), .CK(clk_in), .Q(shmem_addr_i[3]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[113]  ( .D(n868), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[113]) );
  DFF_X1 \shmem_addr_i_reg[2]  ( .D(n194), .CK(clk_in), .Q(shmem_addr_i[2]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[112]  ( .D(n869), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[112]) );
  DFF_X1 \shmem_addr_i_reg[1]  ( .D(n195), .CK(clk_in), .Q(shmem_addr_i[1]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[111]  ( .D(n870), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[111]) );
  DFF_X1 \shmem_addr_i_reg[0]  ( .D(n196), .CK(clk_in), .Q(shmem_addr_i[0]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[110]  ( .D(n871), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[110]) );
  DFF_X1 \warp_id_addr_reg[4]  ( .D(n728), .CK(clk_in), .Q(warp_id_addr[4]), 
        .QN(n267) );
  DFF_X1 \warp_id_addr_reg[3]  ( .D(n727), .CK(clk_in), .Q(warp_id_addr[3]), 
        .QN(n268) );
  DFF_X1 \warp_id_addr_reg[2]  ( .D(n726), .CK(clk_in), .Q(warp_id_addr[2]), 
        .QN(n269) );
  DFF_X1 \warp_id_addr_reg[1]  ( .D(n725), .CK(clk_in), .Q(warp_id_addr[1]), 
        .QN(n270) );
  DFF_X1 \warp_id_addr_reg[0]  ( .D(n724), .CK(clk_in), .Q(warp_id_addr[0]), 
        .QN(n271) );
  DFF_X1 \fence_regs_cta_id_out_reg[25><3]  ( .D(n620), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[25><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[25><2]  ( .D(n621), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[25><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[25><1]  ( .D(n622), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[25><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[25><0]  ( .D(n623), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[25><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[25]  ( .D(n538), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[25]), .QN(n241) );
  DFF_X1 \fence_regs_cta_id_ld_reg[25]  ( .D(n570), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[25]), .QN(n209) );
  DFF_X1 \fence_regs_cta_id_out_reg[17><3]  ( .D(n652), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[17><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[17><2]  ( .D(n653), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[17><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[17><1]  ( .D(n654), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[17><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[17><0]  ( .D(n655), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[17><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[17]  ( .D(n546), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[17]), .QN(n249) );
  DFF_X1 \fence_regs_cta_id_ld_reg[17]  ( .D(n578), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[17]), .QN(n217) );
  DFF_X1 \fence_regs_cta_id_out_reg[9><3]  ( .D(n684), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[9><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[9><2]  ( .D(n685), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[9><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[9><1]  ( .D(n686), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[9><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[9><0]  ( .D(n687), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[9><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[9]  ( .D(n554), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[9]), .QN(n257) );
  DFF_X1 \fence_regs_cta_id_ld_reg[9]  ( .D(n586), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[9]), .QN(n225) );
  DFF_X1 \fence_regs_cta_id_out_reg[1><3]  ( .D(n716), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[1><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[1><2]  ( .D(n717), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[1><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[1><1]  ( .D(n718), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[1><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[1><0]  ( .D(n719), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[1><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[1]  ( .D(n562), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[1]), .QN(n265) );
  DFF_X1 \fence_regs_cta_id_ld_reg[1]  ( .D(n594), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[1]), .QN(n233) );
  DFF_X1 \fence_regs_cta_id_out_reg[27><3]  ( .D(n612), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[27><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[27><2]  ( .D(n613), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[27><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[27><1]  ( .D(n614), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[27><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[27><0]  ( .D(n615), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[27><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[27]  ( .D(n536), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[27]), .QN(n239) );
  DFF_X1 \fence_regs_cta_id_ld_reg[27]  ( .D(n568), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[27]), .QN(n207) );
  DFF_X1 \fence_regs_cta_id_out_reg[19><3]  ( .D(n644), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[19><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[19><2]  ( .D(n645), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[19><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[19><1]  ( .D(n646), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[19><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[19><0]  ( .D(n647), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[19><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[19]  ( .D(n544), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[19]), .QN(n247) );
  DFF_X1 \fence_regs_cta_id_ld_reg[19]  ( .D(n576), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[19]), .QN(n215) );
  DFF_X1 \fence_regs_cta_id_out_reg[11><3]  ( .D(n676), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[11><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[11><2]  ( .D(n677), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[11><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[11><1]  ( .D(n678), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[11><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[11><0]  ( .D(n679), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[11><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[11]  ( .D(n552), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[11]), .QN(n255) );
  DFF_X1 \fence_regs_cta_id_ld_reg[11]  ( .D(n584), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[11]), .QN(n223) );
  DFF_X1 \fence_regs_cta_id_out_reg[3><3]  ( .D(n708), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[3><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[3><2]  ( .D(n709), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[3><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[3><1]  ( .D(n710), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[3><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[3><0]  ( .D(n711), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[3><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[3]  ( .D(n560), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[3]), .QN(n263) );
  DFF_X1 \fence_regs_cta_id_ld_reg[3]  ( .D(n592), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[3]), .QN(n231) );
  DFF_X1 \fence_regs_cta_id_out_reg[29><3]  ( .D(n604), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[29><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[29><2]  ( .D(n605), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[29><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[29><1]  ( .D(n606), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[29><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[29><0]  ( .D(n607), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[29><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[29]  ( .D(n534), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[29]), .QN(n237) );
  DFF_X1 \fence_regs_cta_id_ld_reg[29]  ( .D(n566), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[29]), .QN(n205) );
  DFF_X1 \fence_regs_cta_id_out_reg[21><3]  ( .D(n636), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[21><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[21><2]  ( .D(n637), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[21><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[21><1]  ( .D(n638), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[21><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[21><0]  ( .D(n639), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[21><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[21]  ( .D(n542), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[21]), .QN(n245) );
  DFF_X1 \fence_regs_cta_id_ld_reg[21]  ( .D(n574), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[21]), .QN(n213) );
  DFF_X1 \fence_regs_cta_id_out_reg[13><3]  ( .D(n668), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[13><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[13><2]  ( .D(n669), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[13><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[13><1]  ( .D(n670), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[13><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[13><0]  ( .D(n671), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[13><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[13]  ( .D(n550), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[13]), .QN(n253) );
  DFF_X1 \fence_regs_cta_id_ld_reg[13]  ( .D(n582), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[13]), .QN(n221) );
  DFF_X1 \fence_regs_cta_id_out_reg[5><3]  ( .D(n700), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[5><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[5><2]  ( .D(n701), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[5><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[5><1]  ( .D(n702), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[5><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[5><0]  ( .D(n703), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[5><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[5]  ( .D(n558), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[5]), .QN(n261) );
  DFF_X1 \fence_regs_cta_id_ld_reg[5]  ( .D(n590), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[5]), .QN(n229) );
  DFF_X1 \fence_regs_cta_id_out_reg[31><3]  ( .D(n596), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[31><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[31><2]  ( .D(n597), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[31><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[31><1]  ( .D(n598), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[31><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[31><0]  ( .D(n599), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[31><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[31]  ( .D(n532), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[31]), .QN(n235) );
  DFF_X1 \fence_regs_cta_id_ld_reg[31]  ( .D(n564), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[31]), .QN(n203) );
  DFF_X1 \fence_regs_cta_id_out_reg[23><3]  ( .D(n628), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[23><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[23><2]  ( .D(n629), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[23><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[23><1]  ( .D(n630), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[23><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[23><0]  ( .D(n631), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[23><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[23]  ( .D(n540), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[23]), .QN(n243) );
  DFF_X1 \fence_regs_cta_id_ld_reg[23]  ( .D(n572), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[23]), .QN(n211) );
  DFF_X1 \fence_regs_cta_id_out_reg[15><3]  ( .D(n660), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[15><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[15><2]  ( .D(n661), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[15><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[15><1]  ( .D(n662), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[15><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[15><0]  ( .D(n663), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[15><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[15]  ( .D(n548), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[15]), .QN(n251) );
  DFF_X1 \fence_regs_cta_id_ld_reg[15]  ( .D(n580), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[15]), .QN(n219) );
  DFF_X1 \fence_regs_cta_id_out_reg[7><3]  ( .D(n692), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[7><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[7><2]  ( .D(n693), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[7><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[7><1]  ( .D(n694), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[7><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[7><0]  ( .D(n695), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[7><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[7]  ( .D(n556), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[7]), .QN(n259) );
  DFF_X1 \fence_regs_cta_id_ld_reg[7]  ( .D(n588), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[7]), .QN(n227) );
  DFF_X1 \fence_regs_cta_id_out_reg[24><3]  ( .D(n624), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[24><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[24><2]  ( .D(n625), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[24><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[24><1]  ( .D(n626), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[24><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[24><0]  ( .D(n627), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[24><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[24]  ( .D(n539), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[24]), .QN(n242) );
  DFF_X1 \fence_regs_cta_id_ld_reg[24]  ( .D(n571), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[24]), .QN(n210) );
  DFF_X1 \fence_regs_cta_id_out_reg[16><3]  ( .D(n656), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[16><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[16><2]  ( .D(n657), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[16><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[16><1]  ( .D(n658), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[16><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[16><0]  ( .D(n659), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[16><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[16]  ( .D(n547), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[16]), .QN(n250) );
  DFF_X1 \fence_regs_cta_id_ld_reg[16]  ( .D(n579), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[16]), .QN(n218) );
  DFF_X1 \fence_regs_cta_id_out_reg[8><3]  ( .D(n688), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[8><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[8><2]  ( .D(n689), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[8><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[8><1]  ( .D(n690), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[8><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[8><0]  ( .D(n691), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[8><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[8]  ( .D(n555), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[8]), .QN(n258) );
  DFF_X1 \fence_regs_cta_id_ld_reg[8]  ( .D(n587), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[8]), .QN(n226) );
  DFF_X1 \fence_regs_cta_id_out_reg[0><3]  ( .D(n720), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[0><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[0><2]  ( .D(n721), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[0><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[0><1]  ( .D(n722), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[0><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[0><0]  ( .D(n723), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[0><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[0]  ( .D(n563), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[0]), .QN(n266) );
  DFF_X1 \fence_regs_cta_id_ld_reg[0]  ( .D(n595), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[0]), .QN(n234) );
  DFF_X1 \fence_regs_cta_id_out_reg[26><3]  ( .D(n616), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[26><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[26><2]  ( .D(n617), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[26><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[26><1]  ( .D(n618), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[26><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[26><0]  ( .D(n619), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[26><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[26]  ( .D(n537), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[26]), .QN(n240) );
  DFF_X1 \fence_regs_cta_id_ld_reg[26]  ( .D(n569), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[26]), .QN(n208) );
  DFF_X1 \fence_regs_cta_id_out_reg[18><3]  ( .D(n648), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[18><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[18><2]  ( .D(n649), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[18><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[18><1]  ( .D(n650), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[18><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[18><0]  ( .D(n651), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[18><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[18]  ( .D(n545), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[18]), .QN(n248) );
  DFF_X1 \fence_regs_cta_id_ld_reg[18]  ( .D(n577), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[18]), .QN(n216) );
  DFF_X1 \fence_regs_cta_id_out_reg[10><3]  ( .D(n680), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[10><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[10><2]  ( .D(n681), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[10><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[10><1]  ( .D(n682), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[10><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[10><0]  ( .D(n683), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[10><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[10]  ( .D(n553), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[10]), .QN(n256) );
  DFF_X1 \fence_regs_cta_id_ld_reg[10]  ( .D(n585), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[10]), .QN(n224) );
  DFF_X1 \fence_regs_cta_id_out_reg[2><3]  ( .D(n712), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[2><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[2><2]  ( .D(n713), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[2><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[2><1]  ( .D(n714), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[2><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[2><0]  ( .D(n715), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[2><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[2]  ( .D(n561), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[2]), .QN(n264) );
  DFF_X1 \fence_regs_cta_id_ld_reg[2]  ( .D(n593), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[2]), .QN(n232) );
  DFF_X1 \fence_regs_cta_id_out_reg[28><3]  ( .D(n608), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[28><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[28><2]  ( .D(n609), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[28><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[28><1]  ( .D(n610), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[28><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[28><0]  ( .D(n611), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[28><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[28]  ( .D(n535), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[28]), .QN(n238) );
  DFF_X1 \fence_regs_cta_id_ld_reg[28]  ( .D(n567), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[28]), .QN(n206) );
  DFF_X1 \fence_regs_cta_id_out_reg[20><3]  ( .D(n640), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[20><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[20><2]  ( .D(n641), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[20><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[20><1]  ( .D(n642), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[20><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[20><0]  ( .D(n643), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[20><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[20]  ( .D(n543), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[20]), .QN(n246) );
  DFF_X1 \fence_regs_cta_id_ld_reg[20]  ( .D(n575), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[20]), .QN(n214) );
  DFF_X1 \fence_regs_cta_id_out_reg[12><3]  ( .D(n672), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[12><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[12><2]  ( .D(n673), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[12><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[12><1]  ( .D(n674), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[12><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[12><0]  ( .D(n675), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[12><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[12]  ( .D(n551), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[12]), .QN(n254) );
  DFF_X1 \fence_regs_cta_id_ld_reg[12]  ( .D(n583), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[12]), .QN(n222) );
  DFF_X1 \fence_regs_cta_id_out_reg[4><3]  ( .D(n704), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[4><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[4><2]  ( .D(n705), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[4><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[4><1]  ( .D(n706), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[4><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[4><0]  ( .D(n707), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[4><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[4]  ( .D(n559), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[4]), .QN(n262) );
  DFF_X1 \fence_regs_cta_id_ld_reg[4]  ( .D(n591), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[4]), .QN(n230) );
  DFF_X1 \fence_regs_cta_id_out_reg[30><3]  ( .D(n600), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[30><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[30><2]  ( .D(n601), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[30><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[30><1]  ( .D(n602), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[30><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[30><0]  ( .D(n603), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[30><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[30]  ( .D(n533), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[30]), .QN(n236) );
  DFF_X1 \fence_regs_cta_id_ld_reg[30]  ( .D(n565), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[30]), .QN(n204) );
  DFF_X1 \fence_regs_cta_id_out_reg[22><3]  ( .D(n632), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[22><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[22><2]  ( .D(n633), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[22><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[22><1]  ( .D(n634), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[22><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[22><0]  ( .D(n635), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[22><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[22]  ( .D(n541), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[22]), .QN(n244) );
  DFF_X1 \fence_regs_cta_id_ld_reg[22]  ( .D(n573), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[22]), .QN(n212) );
  DFF_X1 \fence_regs_cta_id_out_reg[14><3]  ( .D(n664), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[14><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[14><2]  ( .D(n665), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[14><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[14><1]  ( .D(n666), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[14><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[14><0]  ( .D(n667), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[14><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[14]  ( .D(n549), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[14]), .QN(n252) );
  DFF_X1 \fence_regs_cta_id_ld_reg[14]  ( .D(n581), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[14]), .QN(n220) );
  DFF_X1 \fence_regs_cta_id_out_reg[6><3]  ( .D(n696), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[6><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[6><2]  ( .D(n697), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[6><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[6><1]  ( .D(n698), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[6><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[6><0]  ( .D(n699), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[6><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[6]  ( .D(n557), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[6]), .QN(n260) );
  DFF_X1 \fence_regs_cta_id_ld_reg[6]  ( .D(n589), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[6]), .QN(n228) );
  NOR2_X2 U313 ( .A1(n439), .A2(n453), .ZN(n438) );
  NOR3_X2 U429 ( .A1(n453), .A2(n496), .A3(n873), .ZN(n495) );
  NAND2_X1 U597 ( .A1(\fence_regs_cta_id_out[31><3] ), .A2(n856), .ZN(n281) );
  NAND2_X1 U598 ( .A1(\fence_regs_cta_id_out[31><2] ), .A2(n856), .ZN(n283) );
  NAND2_X1 U599 ( .A1(\fence_regs_cta_id_out[31><1] ), .A2(n856), .ZN(n285) );
  NAND2_X1 U600 ( .A1(\fence_regs_cta_id_out[31><0] ), .A2(n856), .ZN(n287) );
  NAND2_X1 U601 ( .A1(\fence_regs_cta_id_out[30><3] ), .A2(n855), .ZN(n288) );
  NAND2_X1 U602 ( .A1(\fence_regs_cta_id_out[30><2] ), .A2(n855), .ZN(n289) );
  NAND2_X1 U603 ( .A1(\fence_regs_cta_id_out[30><1] ), .A2(n855), .ZN(n290) );
  NAND2_X1 U604 ( .A1(\fence_regs_cta_id_out[30><0] ), .A2(n855), .ZN(n291) );
  NAND2_X1 U605 ( .A1(\fence_regs_cta_id_out[29><3] ), .A2(n854), .ZN(n292) );
  NAND2_X1 U606 ( .A1(\fence_regs_cta_id_out[29><2] ), .A2(n854), .ZN(n293) );
  NAND2_X1 U607 ( .A1(\fence_regs_cta_id_out[29><1] ), .A2(n854), .ZN(n294) );
  NAND2_X1 U608 ( .A1(\fence_regs_cta_id_out[29><0] ), .A2(n854), .ZN(n295) );
  NAND2_X1 U609 ( .A1(\fence_regs_cta_id_out[28><3] ), .A2(n853), .ZN(n296) );
  NAND2_X1 U610 ( .A1(\fence_regs_cta_id_out[28><2] ), .A2(n853), .ZN(n297) );
  NAND2_X1 U611 ( .A1(\fence_regs_cta_id_out[28><1] ), .A2(n853), .ZN(n298) );
  NAND2_X1 U612 ( .A1(\fence_regs_cta_id_out[28><0] ), .A2(n853), .ZN(n299) );
  NAND2_X1 U613 ( .A1(\fence_regs_cta_id_out[27><3] ), .A2(n852), .ZN(n300) );
  NAND2_X1 U614 ( .A1(\fence_regs_cta_id_out[27><2] ), .A2(n852), .ZN(n301) );
  NAND2_X1 U615 ( .A1(\fence_regs_cta_id_out[27><1] ), .A2(n852), .ZN(n302) );
  NAND2_X1 U616 ( .A1(\fence_regs_cta_id_out[27><0] ), .A2(n852), .ZN(n303) );
  NAND2_X1 U617 ( .A1(\fence_regs_cta_id_out[26><3] ), .A2(n851), .ZN(n304) );
  NAND2_X1 U618 ( .A1(\fence_regs_cta_id_out[26><2] ), .A2(n851), .ZN(n305) );
  NAND2_X1 U619 ( .A1(\fence_regs_cta_id_out[26><1] ), .A2(n851), .ZN(n306) );
  NAND2_X1 U620 ( .A1(\fence_regs_cta_id_out[26><0] ), .A2(n851), .ZN(n307) );
  NAND2_X1 U621 ( .A1(\fence_regs_cta_id_out[25><3] ), .A2(n850), .ZN(n308) );
  NAND2_X1 U622 ( .A1(\fence_regs_cta_id_out[25><2] ), .A2(n850), .ZN(n309) );
  NAND2_X1 U623 ( .A1(\fence_regs_cta_id_out[25><1] ), .A2(n850), .ZN(n310) );
  NAND2_X1 U624 ( .A1(\fence_regs_cta_id_out[25><0] ), .A2(n850), .ZN(n311) );
  NAND2_X1 U625 ( .A1(\fence_regs_cta_id_out[24><3] ), .A2(n849), .ZN(n312) );
  NAND2_X1 U626 ( .A1(\fence_regs_cta_id_out[24><2] ), .A2(n849), .ZN(n313) );
  NAND2_X1 U627 ( .A1(\fence_regs_cta_id_out[24><1] ), .A2(n849), .ZN(n314) );
  NAND2_X1 U628 ( .A1(\fence_regs_cta_id_out[24><0] ), .A2(n849), .ZN(n315) );
  NAND2_X1 U629 ( .A1(\fence_regs_cta_id_out[23><3] ), .A2(n848), .ZN(n316) );
  NAND2_X1 U630 ( .A1(\fence_regs_cta_id_out[23><2] ), .A2(n848), .ZN(n317) );
  NAND2_X1 U631 ( .A1(\fence_regs_cta_id_out[23><1] ), .A2(n848), .ZN(n318) );
  NAND2_X1 U632 ( .A1(\fence_regs_cta_id_out[23><0] ), .A2(n848), .ZN(n319) );
  NAND2_X1 U633 ( .A1(\fence_regs_cta_id_out[22><3] ), .A2(n847), .ZN(n320) );
  NAND2_X1 U634 ( .A1(\fence_regs_cta_id_out[22><2] ), .A2(n847), .ZN(n321) );
  NAND2_X1 U635 ( .A1(\fence_regs_cta_id_out[22><1] ), .A2(n847), .ZN(n322) );
  NAND2_X1 U636 ( .A1(\fence_regs_cta_id_out[22><0] ), .A2(n847), .ZN(n323) );
  NAND2_X1 U637 ( .A1(\fence_regs_cta_id_out[21><3] ), .A2(n846), .ZN(n324) );
  NAND2_X1 U638 ( .A1(\fence_regs_cta_id_out[21><2] ), .A2(n846), .ZN(n325) );
  NAND2_X1 U639 ( .A1(\fence_regs_cta_id_out[21><1] ), .A2(n846), .ZN(n326) );
  NAND2_X1 U640 ( .A1(\fence_regs_cta_id_out[21><0] ), .A2(n846), .ZN(n327) );
  NAND2_X1 U641 ( .A1(\fence_regs_cta_id_out[20><3] ), .A2(n845), .ZN(n328) );
  NAND2_X1 U642 ( .A1(\fence_regs_cta_id_out[20><2] ), .A2(n845), .ZN(n329) );
  NAND2_X1 U643 ( .A1(\fence_regs_cta_id_out[20><1] ), .A2(n845), .ZN(n330) );
  NAND2_X1 U644 ( .A1(\fence_regs_cta_id_out[20><0] ), .A2(n845), .ZN(n331) );
  NAND2_X1 U645 ( .A1(\fence_regs_cta_id_out[19><3] ), .A2(n844), .ZN(n332) );
  NAND2_X1 U646 ( .A1(\fence_regs_cta_id_out[19><2] ), .A2(n844), .ZN(n333) );
  NAND2_X1 U647 ( .A1(\fence_regs_cta_id_out[19><1] ), .A2(n844), .ZN(n334) );
  NAND2_X1 U648 ( .A1(\fence_regs_cta_id_out[19><0] ), .A2(n844), .ZN(n335) );
  NAND2_X1 U649 ( .A1(\fence_regs_cta_id_out[18><3] ), .A2(n843), .ZN(n336) );
  NAND2_X1 U650 ( .A1(\fence_regs_cta_id_out[18><2] ), .A2(n843), .ZN(n337) );
  NAND2_X1 U651 ( .A1(\fence_regs_cta_id_out[18><1] ), .A2(n843), .ZN(n338) );
  NAND2_X1 U652 ( .A1(\fence_regs_cta_id_out[18><0] ), .A2(n843), .ZN(n339) );
  NAND2_X1 U653 ( .A1(\fence_regs_cta_id_out[17><3] ), .A2(n842), .ZN(n340) );
  NAND2_X1 U654 ( .A1(\fence_regs_cta_id_out[17><2] ), .A2(n842), .ZN(n341) );
  NAND2_X1 U655 ( .A1(\fence_regs_cta_id_out[17><1] ), .A2(n842), .ZN(n342) );
  NAND2_X1 U656 ( .A1(\fence_regs_cta_id_out[17><0] ), .A2(n842), .ZN(n343) );
  NAND2_X1 U657 ( .A1(\fence_regs_cta_id_out[16><3] ), .A2(n841), .ZN(n344) );
  NAND2_X1 U658 ( .A1(\fence_regs_cta_id_out[16><2] ), .A2(n841), .ZN(n345) );
  NAND2_X1 U659 ( .A1(\fence_regs_cta_id_out[16><1] ), .A2(n841), .ZN(n346) );
  NAND2_X1 U660 ( .A1(\fence_regs_cta_id_out[16><0] ), .A2(n841), .ZN(n347) );
  NAND2_X1 U661 ( .A1(\fence_regs_cta_id_out[15><3] ), .A2(n840), .ZN(n348) );
  NAND2_X1 U662 ( .A1(\fence_regs_cta_id_out[15><2] ), .A2(n840), .ZN(n349) );
  NAND2_X1 U663 ( .A1(\fence_regs_cta_id_out[15><1] ), .A2(n840), .ZN(n350) );
  NAND2_X1 U664 ( .A1(\fence_regs_cta_id_out[15><0] ), .A2(n840), .ZN(n351) );
  NAND2_X1 U665 ( .A1(\fence_regs_cta_id_out[14><3] ), .A2(n839), .ZN(n352) );
  NAND2_X1 U666 ( .A1(\fence_regs_cta_id_out[14><2] ), .A2(n839), .ZN(n353) );
  NAND2_X1 U667 ( .A1(\fence_regs_cta_id_out[14><1] ), .A2(n839), .ZN(n354) );
  NAND2_X1 U668 ( .A1(\fence_regs_cta_id_out[14><0] ), .A2(n839), .ZN(n355) );
  NAND2_X1 U669 ( .A1(\fence_regs_cta_id_out[13><3] ), .A2(n838), .ZN(n356) );
  NAND2_X1 U670 ( .A1(\fence_regs_cta_id_out[13><2] ), .A2(n838), .ZN(n357) );
  NAND2_X1 U671 ( .A1(\fence_regs_cta_id_out[13><1] ), .A2(n838), .ZN(n358) );
  NAND2_X1 U672 ( .A1(\fence_regs_cta_id_out[13><0] ), .A2(n838), .ZN(n359) );
  NAND2_X1 U673 ( .A1(\fence_regs_cta_id_out[12><3] ), .A2(n837), .ZN(n360) );
  NAND2_X1 U674 ( .A1(\fence_regs_cta_id_out[12><2] ), .A2(n837), .ZN(n361) );
  NAND2_X1 U675 ( .A1(\fence_regs_cta_id_out[12><1] ), .A2(n837), .ZN(n362) );
  NAND2_X1 U676 ( .A1(\fence_regs_cta_id_out[12><0] ), .A2(n837), .ZN(n363) );
  NAND2_X1 U677 ( .A1(\fence_regs_cta_id_out[11><3] ), .A2(n836), .ZN(n364) );
  NAND2_X1 U678 ( .A1(\fence_regs_cta_id_out[11><2] ), .A2(n836), .ZN(n365) );
  NAND2_X1 U679 ( .A1(\fence_regs_cta_id_out[11><1] ), .A2(n836), .ZN(n366) );
  NAND2_X1 U680 ( .A1(\fence_regs_cta_id_out[11><0] ), .A2(n836), .ZN(n367) );
  NAND2_X1 U681 ( .A1(\fence_regs_cta_id_out[10><3] ), .A2(n835), .ZN(n368) );
  NAND2_X1 U682 ( .A1(\fence_regs_cta_id_out[10><2] ), .A2(n835), .ZN(n369) );
  NAND2_X1 U683 ( .A1(\fence_regs_cta_id_out[10><1] ), .A2(n835), .ZN(n370) );
  NAND2_X1 U684 ( .A1(\fence_regs_cta_id_out[10><0] ), .A2(n835), .ZN(n371) );
  NAND2_X1 U685 ( .A1(\fence_regs_cta_id_out[9><3] ), .A2(n834), .ZN(n372) );
  NAND2_X1 U686 ( .A1(\fence_regs_cta_id_out[9><2] ), .A2(n834), .ZN(n373) );
  NAND2_X1 U687 ( .A1(\fence_regs_cta_id_out[9><1] ), .A2(n834), .ZN(n374) );
  NAND2_X1 U688 ( .A1(\fence_regs_cta_id_out[9><0] ), .A2(n834), .ZN(n375) );
  NAND2_X1 U689 ( .A1(\fence_regs_cta_id_out[8><3] ), .A2(n833), .ZN(n376) );
  NAND2_X1 U690 ( .A1(\fence_regs_cta_id_out[8><2] ), .A2(n833), .ZN(n377) );
  NAND2_X1 U691 ( .A1(\fence_regs_cta_id_out[8><1] ), .A2(n833), .ZN(n378) );
  NAND2_X1 U692 ( .A1(\fence_regs_cta_id_out[8><0] ), .A2(n833), .ZN(n379) );
  NAND2_X1 U693 ( .A1(\fence_regs_cta_id_out[7><3] ), .A2(n832), .ZN(n380) );
  NAND2_X1 U694 ( .A1(\fence_regs_cta_id_out[7><2] ), .A2(n832), .ZN(n381) );
  NAND2_X1 U695 ( .A1(\fence_regs_cta_id_out[7><1] ), .A2(n832), .ZN(n382) );
  NAND2_X1 U696 ( .A1(\fence_regs_cta_id_out[7><0] ), .A2(n832), .ZN(n383) );
  NAND2_X1 U697 ( .A1(\fence_regs_cta_id_out[6><3] ), .A2(n831), .ZN(n384) );
  NAND2_X1 U698 ( .A1(\fence_regs_cta_id_out[6><2] ), .A2(n831), .ZN(n385) );
  NAND2_X1 U699 ( .A1(\fence_regs_cta_id_out[6><1] ), .A2(n831), .ZN(n386) );
  NAND2_X1 U700 ( .A1(\fence_regs_cta_id_out[6><0] ), .A2(n831), .ZN(n387) );
  NAND2_X1 U701 ( .A1(\fence_regs_cta_id_out[5><3] ), .A2(n830), .ZN(n388) );
  NAND2_X1 U702 ( .A1(\fence_regs_cta_id_out[5><2] ), .A2(n830), .ZN(n389) );
  NAND2_X1 U703 ( .A1(\fence_regs_cta_id_out[5><1] ), .A2(n830), .ZN(n390) );
  NAND2_X1 U704 ( .A1(\fence_regs_cta_id_out[5><0] ), .A2(n830), .ZN(n391) );
  NAND2_X1 U705 ( .A1(\fence_regs_cta_id_out[4><3] ), .A2(n829), .ZN(n392) );
  NAND2_X1 U706 ( .A1(\fence_regs_cta_id_out[4><2] ), .A2(n829), .ZN(n393) );
  NAND2_X1 U707 ( .A1(\fence_regs_cta_id_out[4><1] ), .A2(n829), .ZN(n394) );
  NAND2_X1 U708 ( .A1(\fence_regs_cta_id_out[4><0] ), .A2(n829), .ZN(n395) );
  NAND2_X1 U709 ( .A1(\fence_regs_cta_id_out[3><3] ), .A2(n828), .ZN(n396) );
  NAND2_X1 U710 ( .A1(\fence_regs_cta_id_out[3><2] ), .A2(n828), .ZN(n397) );
  NAND2_X1 U711 ( .A1(\fence_regs_cta_id_out[3><1] ), .A2(n828), .ZN(n398) );
  NAND2_X1 U712 ( .A1(\fence_regs_cta_id_out[3><0] ), .A2(n828), .ZN(n399) );
  NAND2_X1 U713 ( .A1(\fence_regs_cta_id_out[2><3] ), .A2(n827), .ZN(n400) );
  NAND2_X1 U714 ( .A1(\fence_regs_cta_id_out[2><2] ), .A2(n827), .ZN(n401) );
  NAND2_X1 U715 ( .A1(\fence_regs_cta_id_out[2><1] ), .A2(n827), .ZN(n402) );
  NAND2_X1 U716 ( .A1(\fence_regs_cta_id_out[2><0] ), .A2(n827), .ZN(n403) );
  NAND2_X1 U717 ( .A1(\fence_regs_cta_id_out[1><3] ), .A2(n826), .ZN(n404) );
  NAND2_X1 U718 ( .A1(\fence_regs_cta_id_out[1><2] ), .A2(n826), .ZN(n405) );
  NAND2_X1 U719 ( .A1(\fence_regs_cta_id_out[1><1] ), .A2(n826), .ZN(n406) );
  NAND2_X1 U720 ( .A1(\fence_regs_cta_id_out[1><0] ), .A2(n826), .ZN(n407) );
  NAND2_X1 U721 ( .A1(\fence_regs_cta_id_out[0><3] ), .A2(n825), .ZN(n408) );
  NAND2_X1 U722 ( .A1(block_num_i[3]), .A2(n34), .ZN(n280) );
  NAND2_X1 U723 ( .A1(\fence_regs_cta_id_out[0><2] ), .A2(n825), .ZN(n409) );
  NAND2_X1 U724 ( .A1(block_num_i[2]), .A2(n34), .ZN(n282) );
  NAND2_X1 U725 ( .A1(\fence_regs_cta_id_out[0><1] ), .A2(n825), .ZN(n410) );
  NAND2_X1 U726 ( .A1(block_num_i[1]), .A2(n35), .ZN(n284) );
  NAND2_X1 U727 ( .A1(\fence_regs_cta_id_out[0><0] ), .A2(n825), .ZN(n411) );
  NAND2_X1 U728 ( .A1(block_num_i[0]), .A2(n35), .ZN(n286) );
  NAND2_X1 U731 ( .A1(n455), .A2(n460), .ZN(n797) );
  NAND2_X1 U732 ( .A1(warp_gen_done), .A2(n461), .ZN(n460) );
  NAND2_X1 U733 ( .A1(warp_num_i[0]), .A2(n475), .ZN(n474) );
  NAND2_X1 U734 ( .A1(warp_num_i[1]), .A2(n475), .ZN(n476) );
  NAND2_X1 U735 ( .A1(warp_num_i[2]), .A2(n475), .ZN(n477) );
  NAND2_X1 U736 ( .A1(warp_num_i[3]), .A2(n475), .ZN(n478) );
  NAND2_X1 U737 ( .A1(warp_num_i[4]), .A2(n475), .ZN(n479) );
  NAND2_X1 U738 ( .A1(n872), .A2(n274), .ZN(n473) );
  NAND2_X1 U739 ( .A1(block_num_cnt[1]), .A2(n142), .ZN(n485) );
  NAND3_X1 U740 ( .A1(n275), .A2(n145), .A3(n872), .ZN(n487) );
  NAND3_X1 U741 ( .A1(n872), .A2(n275), .A3(block_num_cnt[0]), .ZN(n483) );
  NAND2_X1 U742 ( .A1(n489), .A2(n22), .ZN(n812) );
  NAND2_X1 U743 ( .A1(warp_state_wr_en_out), .A2(n490), .ZN(n489) );
  NAND2_X1 U744 ( .A1(n491), .A2(n22), .ZN(n813) );
  NAND2_X1 U745 ( .A1(warp_pool_wr_en_out), .A2(n490), .ZN(n491) );
  NAND3_X1 U746 ( .A1(n202), .A2(n201), .A3(warp_generator_state_machine[2]), 
        .ZN(n455) );
  NAND3_X1 U747 ( .A1(warp_id_addr[3]), .A2(n528), .A3(warp_id_addr[4]), .ZN(
        n518) );
  NAND3_X1 U748 ( .A1(n528), .A2(n268), .A3(warp_id_addr[4]), .ZN(n529) );
  NAND3_X1 U749 ( .A1(n528), .A2(n267), .A3(warp_id_addr[3]), .ZN(n530) );
  NAND3_X1 U750 ( .A1(warp_id_addr[1]), .A2(warp_id_addr[0]), .A3(
        warp_id_addr[2]), .ZN(n519) );
  NAND3_X1 U751 ( .A1(warp_id_addr[1]), .A2(n271), .A3(warp_id_addr[2]), .ZN(
        n521) );
  NAND3_X1 U752 ( .A1(warp_id_addr[0]), .A2(n270), .A3(warp_id_addr[2]), .ZN(
        n522) );
  NAND3_X1 U753 ( .A1(n271), .A2(n270), .A3(warp_id_addr[2]), .ZN(n523) );
  NAND3_X1 U754 ( .A1(warp_id_addr[0]), .A2(n269), .A3(warp_id_addr[1]), .ZN(
        n524) );
  NAND3_X1 U755 ( .A1(n271), .A2(n269), .A3(warp_id_addr[1]), .ZN(n525) );
  NAND3_X1 U756 ( .A1(n270), .A2(n269), .A3(warp_id_addr[0]), .ZN(n526) );
  NAND3_X1 U757 ( .A1(n201), .A2(n200), .A3(warp_generator_state_machine[0]), 
        .ZN(n453) );
  NAND3_X1 U758 ( .A1(n268), .A2(n267), .A3(n528), .ZN(n531) );
  NAND3_X1 U759 ( .A1(n270), .A2(n269), .A3(n271), .ZN(n527) );
  NAND3_X1 U762 ( .A1(n201), .A2(n200), .A3(n202), .ZN(n461) );
  warp_id_calc uWarpIdCalc ( .clk(clk_in), .reset(n119), .en(
        warp_id_calc_en_i), .block_num_in(block_num_i), .gprs_size_in(
        gprs_size_in), .warp_num_in(warp_num_i), .warps_per_block_in(
        warps_per_block_in), .gprs_base_addr_out(gprs_base_addr_o), 
        .warp_id_out(warp_id_o) );
  warp_generator_SHMEM_ADDR_SIZE14_DW01_inc_1 add_127 ( .A(warps_per_block_cnt), .SUM({N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92}) );
  warp_generator_SHMEM_ADDR_SIZE14_DW02_mult_0 mult_124 ( .A(block_num_cnt), 
        .B(shmem_size_in[13:0]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, N77, N76, N75, N74, N73, N72, N71, N70, N69, 
        N68, N67, N66, N65, N64}) );
  warp_generator_SHMEM_ADDR_SIZE14_DW01_add_0 add_124 ( .A(
        shmem_base_addr_in[13:0]), .B({N77, N76, N75, N74, N73, N72, N71, N70, 
        N69, N68, N67, N66, N65, N64}), .CI(1'b0), .SUM({N91, N90, N89, N88, 
        N87, N86, N85, N84, N83, N82, N81, N80, N79, N78}) );
  HA_X1 \add_155/U1_1_1  ( .A(warp_id_o[1]), .B(warp_id_o[0]), .CO(
        \add_155/carry[2] ), .S(N254) );
  HA_X1 \add_155/U1_1_2  ( .A(warp_id_o[2]), .B(\add_155/carry[2] ), .CO(
        \add_155/carry[3] ), .S(N255) );
  HA_X1 \add_155/U1_1_3  ( .A(warp_id_o[3]), .B(\add_155/carry[3] ), .CO(
        \add_155/carry[4] ), .S(N256) );
  INV_X1 U11 ( .A(n133), .ZN(n139) );
  NOR3_X1 U75 ( .A1(warp_generator_state_machine[0]), .A2(
        warp_generator_state_machine[2]), .A3(n201), .ZN(n413) );
  AND3_X1 U76 ( .A1(warp_generator_state_machine[0]), .A2(n200), .A3(
        warp_generator_state_machine[1]), .ZN(n1) );
  AND2_X1 U77 ( .A1(n461), .A2(n24), .ZN(n3) );
  INV_X1 U78 ( .A(n49), .ZN(n38) );
  INV_X1 U79 ( .A(n48), .ZN(n37) );
  INV_X1 U80 ( .A(n47), .ZN(n36) );
  NAND2_X1 U81 ( .A1(n274), .A2(n126), .ZN(n439) );
  BUF_X1 U82 ( .A(n52), .Z(n50) );
  BUF_X1 U83 ( .A(n52), .Z(n49) );
  BUF_X1 U84 ( .A(n117), .Z(n48) );
  BUF_X1 U85 ( .A(n117), .Z(n47) );
  BUF_X1 U86 ( .A(n117), .Z(n46) );
  INV_X1 U87 ( .A(n488), .ZN(n275) );
  BUF_X1 U88 ( .A(n520), .Z(n4) );
  BUF_X1 U89 ( .A(n520), .Z(n5) );
  BUF_X1 U90 ( .A(n520), .Z(n6) );
  BUF_X1 U91 ( .A(n118), .Z(n39) );
  BUF_X1 U92 ( .A(n118), .Z(n44) );
  BUF_X1 U93 ( .A(n118), .Z(n45) );
  BUF_X1 U94 ( .A(n52), .Z(n51) );
  NOR2_X2 U95 ( .A1(n857), .A2(n480), .ZN(n496) );
  INV_X1 U96 ( .A(N869), .ZN(n831) );
  INV_X1 U97 ( .A(N877), .ZN(n839) );
  INV_X1 U98 ( .A(N885), .ZN(n847) );
  INV_X1 U99 ( .A(N867), .ZN(n829) );
  INV_X1 U100 ( .A(N875), .ZN(n837) );
  INV_X1 U101 ( .A(N883), .ZN(n845) );
  INV_X1 U102 ( .A(N865), .ZN(n827) );
  INV_X1 U103 ( .A(N873), .ZN(n835) );
  INV_X1 U104 ( .A(N881), .ZN(n843) );
  INV_X1 U105 ( .A(N863), .ZN(n825) );
  INV_X1 U106 ( .A(N871), .ZN(n833) );
  INV_X1 U107 ( .A(N879), .ZN(n841) );
  INV_X1 U108 ( .A(N870), .ZN(n832) );
  INV_X1 U109 ( .A(N878), .ZN(n840) );
  INV_X1 U110 ( .A(N886), .ZN(n848) );
  INV_X1 U111 ( .A(N868), .ZN(n830) );
  INV_X1 U112 ( .A(N876), .ZN(n838) );
  INV_X1 U113 ( .A(N884), .ZN(n846) );
  INV_X1 U114 ( .A(N866), .ZN(n828) );
  INV_X1 U115 ( .A(N874), .ZN(n836) );
  INV_X1 U116 ( .A(N882), .ZN(n844) );
  INV_X1 U117 ( .A(N864), .ZN(n826) );
  INV_X1 U118 ( .A(N872), .ZN(n834) );
  INV_X1 U119 ( .A(N880), .ZN(n842) );
  INV_X1 U120 ( .A(N893), .ZN(n855) );
  INV_X1 U121 ( .A(N891), .ZN(n853) );
  INV_X1 U122 ( .A(N889), .ZN(n851) );
  INV_X1 U123 ( .A(N887), .ZN(n849) );
  INV_X1 U124 ( .A(N894), .ZN(n856) );
  INV_X1 U125 ( .A(N892), .ZN(n854) );
  INV_X1 U126 ( .A(N890), .ZN(n852) );
  INV_X1 U127 ( .A(N888), .ZN(n850) );
  INV_X1 U128 ( .A(n475), .ZN(n274) );
  AOI21_X1 U129 ( .B1(n873), .B2(n480), .A(n857), .ZN(n488) );
  NOR2_X1 U130 ( .A1(n23), .A2(n119), .ZN(n528) );
  NOR2_X1 U131 ( .A1(n872), .A2(n38), .ZN(n490) );
  BUF_X1 U132 ( .A(n3), .Z(n52) );
  BUF_X1 U133 ( .A(n3), .Z(n117) );
  INV_X1 U134 ( .A(n34), .ZN(n24) );
  INV_X1 U135 ( .A(n33), .ZN(n22) );
  INV_X1 U136 ( .A(n33), .ZN(n21) );
  INV_X1 U137 ( .A(n31), .ZN(n20) );
  INV_X1 U138 ( .A(n30), .ZN(n19) );
  INV_X1 U139 ( .A(n412), .ZN(n199) );
  OAI21_X1 U140 ( .B1(n872), .B2(n857), .A(n121), .ZN(n520) );
  BUF_X1 U141 ( .A(n3), .Z(n118) );
  INV_X1 U142 ( .A(n119), .ZN(n121) );
  NOR2_X1 U143 ( .A1(n453), .A2(n508), .ZN(n480) );
  AOI21_X1 U144 ( .B1(n480), .B2(N62), .A(n857), .ZN(n475) );
  OAI21_X1 U145 ( .B1(n518), .B2(n521), .A(n6), .ZN(N893) );
  OAI21_X1 U146 ( .B1(n518), .B2(n523), .A(n6), .ZN(N891) );
  OAI21_X1 U147 ( .B1(n518), .B2(n525), .A(n6), .ZN(N889) );
  OAI21_X1 U148 ( .B1(n518), .B2(n527), .A(n6), .ZN(N887) );
  OAI21_X1 U149 ( .B1(n518), .B2(n519), .A(n6), .ZN(N894) );
  OAI21_X1 U150 ( .B1(n518), .B2(n522), .A(n6), .ZN(N892) );
  OAI21_X1 U151 ( .B1(n518), .B2(n524), .A(n6), .ZN(N890) );
  OAI21_X1 U152 ( .B1(n518), .B2(n526), .A(n6), .ZN(N888) );
  OAI21_X1 U153 ( .B1(n521), .B2(n531), .A(n4), .ZN(N869) );
  OAI21_X1 U154 ( .B1(n523), .B2(n531), .A(n4), .ZN(N867) );
  OAI21_X1 U155 ( .B1(n525), .B2(n531), .A(n4), .ZN(N865) );
  OAI21_X1 U156 ( .B1(n527), .B2(n531), .A(n4), .ZN(N863) );
  OAI21_X1 U157 ( .B1(n519), .B2(n531), .A(n4), .ZN(N870) );
  OAI21_X1 U158 ( .B1(n522), .B2(n531), .A(n4), .ZN(N868) );
  OAI21_X1 U159 ( .B1(n524), .B2(n531), .A(n4), .ZN(N866) );
  OAI21_X1 U160 ( .B1(n526), .B2(n531), .A(n4), .ZN(N864) );
  OAI21_X1 U161 ( .B1(n521), .B2(n530), .A(n5), .ZN(N877) );
  OAI21_X1 U162 ( .B1(n521), .B2(n529), .A(n5), .ZN(N885) );
  OAI21_X1 U163 ( .B1(n523), .B2(n530), .A(n5), .ZN(N875) );
  OAI21_X1 U164 ( .B1(n523), .B2(n529), .A(n5), .ZN(N883) );
  OAI21_X1 U165 ( .B1(n525), .B2(n530), .A(n4), .ZN(N873) );
  OAI21_X1 U166 ( .B1(n525), .B2(n529), .A(n5), .ZN(N881) );
  OAI21_X1 U167 ( .B1(n527), .B2(n530), .A(n4), .ZN(N871) );
  OAI21_X1 U168 ( .B1(n527), .B2(n529), .A(n5), .ZN(N879) );
  OAI21_X1 U169 ( .B1(n519), .B2(n530), .A(n5), .ZN(N878) );
  OAI21_X1 U170 ( .B1(n519), .B2(n529), .A(n5), .ZN(N886) );
  OAI21_X1 U171 ( .B1(n522), .B2(n530), .A(n5), .ZN(N876) );
  OAI21_X1 U172 ( .B1(n522), .B2(n529), .A(n5), .ZN(N884) );
  OAI21_X1 U173 ( .B1(n524), .B2(n530), .A(n4), .ZN(N874) );
  OAI21_X1 U174 ( .B1(n524), .B2(n529), .A(n5), .ZN(N882) );
  OAI21_X1 U175 ( .B1(n526), .B2(n530), .A(n4), .ZN(N872) );
  OAI21_X1 U176 ( .B1(n526), .B2(n529), .A(n5), .ZN(N880) );
  INV_X1 U177 ( .A(N62), .ZN(n873) );
  BUF_X1 U178 ( .A(n1), .Z(n34) );
  BUF_X1 U179 ( .A(n1), .Z(n33) );
  INV_X1 U180 ( .A(n492), .ZN(n198) );
  INV_X1 U181 ( .A(n453), .ZN(n872) );
  BUF_X1 U182 ( .A(n282), .Z(n13) );
  BUF_X1 U183 ( .A(n280), .Z(n16) );
  BUF_X1 U184 ( .A(n282), .Z(n14) );
  BUF_X1 U185 ( .A(n280), .Z(n17) );
  BUF_X1 U186 ( .A(n286), .Z(n7) );
  BUF_X1 U187 ( .A(n284), .Z(n10) );
  BUF_X1 U188 ( .A(n286), .Z(n8) );
  BUF_X1 U189 ( .A(n284), .Z(n11) );
  INV_X1 U190 ( .A(n455), .ZN(n272) );
  INV_X1 U191 ( .A(n461), .ZN(n857) );
  BUF_X1 U192 ( .A(n282), .Z(n15) );
  BUF_X1 U193 ( .A(n280), .Z(n18) );
  BUF_X1 U194 ( .A(n286), .Z(n9) );
  BUF_X1 U195 ( .A(n284), .Z(n12) );
  BUF_X1 U196 ( .A(n1), .Z(n28) );
  BUF_X1 U197 ( .A(n1), .Z(n29) );
  BUF_X1 U198 ( .A(n1), .Z(n30) );
  BUF_X1 U199 ( .A(n1), .Z(n32) );
  BUF_X1 U200 ( .A(n1), .Z(n31) );
  BUF_X1 U201 ( .A(n1), .Z(n25) );
  BUF_X1 U202 ( .A(n1), .Z(n26) );
  BUF_X1 U203 ( .A(n1), .Z(n27) );
  BUF_X1 U204 ( .A(n1), .Z(n35) );
  BUF_X1 U205 ( .A(host_reset), .Z(n119) );
  BUF_X1 U206 ( .A(host_reset), .Z(n120) );
  INV_X1 U207 ( .A(n458), .ZN(n162) );
  AOI22_X1 U208 ( .A1(N257), .A2(n272), .B1(num_warps_out[4]), .B2(n455), .ZN(
        n458) );
  INV_X1 U209 ( .A(n456), .ZN(n170) );
  AOI22_X1 U210 ( .A1(N255), .A2(n272), .B1(num_warps_out[2]), .B2(n455), .ZN(
        n456) );
  INV_X1 U211 ( .A(n452), .ZN(n183) );
  AOI22_X1 U212 ( .A1(N91), .A2(n438), .B1(shmem_addr_i[13]), .B2(n439), .ZN(
        n452) );
  INV_X1 U213 ( .A(n454), .ZN(n174) );
  AOI22_X1 U214 ( .A1(N254), .A2(n272), .B1(num_warps_out[1]), .B2(n455), .ZN(
        n454) );
  INV_X1 U215 ( .A(n457), .ZN(n166) );
  AOI22_X1 U216 ( .A1(N256), .A2(n272), .B1(num_warps_out[3]), .B2(n455), .ZN(
        n457) );
  INV_X1 U217 ( .A(n468), .ZN(n168) );
  AOI22_X1 U218 ( .A1(n50), .A2(warp_pool_addr_out[3]), .B1(n32), .B2(
        warp_id_o[3]), .ZN(n468) );
  INV_X1 U219 ( .A(n463), .ZN(n169) );
  AOI22_X1 U220 ( .A1(n49), .A2(warp_state_addr_out[3]), .B1(n31), .B2(
        warp_id_o[3]), .ZN(n463) );
  INV_X1 U221 ( .A(n469), .ZN(n172) );
  AOI22_X1 U222 ( .A1(n50), .A2(warp_pool_addr_out[2]), .B1(n32), .B2(
        warp_id_o[2]), .ZN(n469) );
  INV_X1 U223 ( .A(n464), .ZN(n173) );
  AOI22_X1 U224 ( .A1(n49), .A2(warp_state_addr_out[2]), .B1(n31), .B2(
        warp_id_o[2]), .ZN(n464) );
  INV_X1 U225 ( .A(n470), .ZN(n176) );
  AOI22_X1 U226 ( .A1(n50), .A2(warp_pool_addr_out[1]), .B1(n32), .B2(
        warp_id_o[1]), .ZN(n470) );
  INV_X1 U227 ( .A(n465), .ZN(n177) );
  AOI22_X1 U228 ( .A1(n49), .A2(warp_state_addr_out[1]), .B1(n31), .B2(
        warp_id_o[1]), .ZN(n465) );
  INV_X1 U229 ( .A(n467), .ZN(n164) );
  AOI22_X1 U230 ( .A1(n50), .A2(warp_pool_addr_out[4]), .B1(n32), .B2(
        warp_id_o[4]), .ZN(n467) );
  INV_X1 U231 ( .A(n462), .ZN(n165) );
  AOI22_X1 U232 ( .A1(n48), .A2(warp_state_addr_out[4]), .B1(n30), .B2(
        warp_id_o[4]), .ZN(n462) );
  INV_X1 U233 ( .A(warps_per_block_in[4]), .ZN(n137) );
  INV_X1 U234 ( .A(n502), .ZN(n818) );
  AOI22_X1 U235 ( .A1(warps_per_block_cnt[4]), .A2(n496), .B1(n495), .B2(N96), 
        .ZN(n502) );
  INV_X1 U236 ( .A(n503), .ZN(n817) );
  AOI22_X1 U237 ( .A1(warps_per_block_cnt[3]), .A2(n496), .B1(n495), .B2(N95), 
        .ZN(n503) );
  INV_X1 U238 ( .A(n504), .ZN(n816) );
  AOI22_X1 U239 ( .A1(warps_per_block_cnt[2]), .A2(n496), .B1(n495), .B2(N94), 
        .ZN(n504) );
  INV_X1 U240 ( .A(n505), .ZN(n279) );
  AOI22_X1 U241 ( .A1(warps_per_block_cnt[1]), .A2(n496), .B1(n495), .B2(N93), 
        .ZN(n505) );
  INV_X1 U242 ( .A(n506), .ZN(n278) );
  AOI22_X1 U243 ( .A1(warps_per_block_cnt[0]), .A2(n496), .B1(n495), .B2(N92), 
        .ZN(n506) );
  NAND4_X1 U244 ( .A1(n455), .A2(n19), .A3(n511), .A4(n512), .ZN(n492) );
  AOI21_X1 U245 ( .B1(en), .B2(n857), .A(n413), .ZN(n512) );
  OAI21_X1 U246 ( .B1(n508), .B2(N62), .A(n872), .ZN(n511) );
  INV_X1 U247 ( .A(n130), .ZN(n138) );
  AOI21_X1 U248 ( .B1(n141), .B2(num_blocks_in[3]), .A(n874), .ZN(n508) );
  INV_X1 U249 ( .A(n513), .ZN(n874) );
  OAI222_X1 U250 ( .A1(n875), .A2(n142), .B1(num_blocks_in[2]), .B2(n514), 
        .C1(num_blocks_in[3]), .C2(n141), .ZN(n513) );
  INV_X1 U251 ( .A(n515), .ZN(n875) );
  OAI21_X1 U252 ( .B1(block_num_cnt[1]), .B2(n453), .A(n486), .ZN(n484) );
  AOI21_X1 U253 ( .B1(n145), .B2(n872), .A(n488), .ZN(n486) );
  OAI22_X1 U254 ( .A1(n155), .A2(n274), .B1(n473), .B2(n145), .ZN(n807) );
  OAI21_X1 U255 ( .B1(n516), .B2(num_blocks_in[1]), .A(n517), .ZN(n515) );
  OAI21_X1 U256 ( .B1(block_num_cnt[0]), .B2(n876), .A(block_num_cnt[1]), .ZN(
        n517) );
  NOR3_X1 U257 ( .A1(n876), .A2(block_num_cnt[1]), .A3(block_num_cnt[0]), .ZN(
        n516) );
  INV_X1 U258 ( .A(num_blocks_in[0]), .ZN(n876) );
  OAI22_X1 U259 ( .A1(n152), .A2(n274), .B1(n141), .B2(n473), .ZN(n801) );
  OAI22_X1 U260 ( .A1(n153), .A2(n274), .B1(n142), .B2(n473), .ZN(n800) );
  OAI22_X1 U261 ( .A1(n154), .A2(n274), .B1(n143), .B2(n473), .ZN(n799) );
  OAI22_X1 U262 ( .A1(n412), .A2(n175), .B1(n199), .B2(n270), .ZN(n725) );
  INV_X1 U263 ( .A(warp_id_o[1]), .ZN(n175) );
  OAI22_X1 U264 ( .A1(n412), .A2(n171), .B1(n199), .B2(n269), .ZN(n726) );
  INV_X1 U265 ( .A(warp_id_o[2]), .ZN(n171) );
  OAI22_X1 U266 ( .A1(n412), .A2(n167), .B1(n199), .B2(n268), .ZN(n727) );
  INV_X1 U267 ( .A(warp_id_o[3]), .ZN(n167) );
  OAI22_X1 U268 ( .A1(n412), .A2(n163), .B1(n199), .B2(n267), .ZN(n728) );
  INV_X1 U269 ( .A(warp_id_o[4]), .ZN(n163) );
  OAI22_X1 U270 ( .A1(n276), .A2(n142), .B1(n483), .B2(n485), .ZN(n809) );
  INV_X1 U271 ( .A(n484), .ZN(n276) );
  OAI22_X1 U272 ( .A1(n839), .A2(n21), .B1(N877), .B2(n220), .ZN(n581) );
  OAI22_X1 U273 ( .A1(n839), .A2(n21), .B1(N877), .B2(n252), .ZN(n549) );
  OAI22_X1 U274 ( .A1(n847), .A2(n19), .B1(N885), .B2(n212), .ZN(n573) );
  OAI22_X1 U275 ( .A1(n847), .A2(n22), .B1(N885), .B2(n244), .ZN(n541) );
  OAI22_X1 U276 ( .A1(n837), .A2(n21), .B1(N875), .B2(n222), .ZN(n583) );
  OAI22_X1 U277 ( .A1(n837), .A2(n19), .B1(N875), .B2(n254), .ZN(n551) );
  OAI22_X1 U278 ( .A1(n845), .A2(n20), .B1(N883), .B2(n214), .ZN(n575) );
  OAI22_X1 U279 ( .A1(n845), .A2(n20), .B1(N883), .B2(n246), .ZN(n543) );
  OAI22_X1 U280 ( .A1(n835), .A2(n21), .B1(N873), .B2(n224), .ZN(n585) );
  OAI22_X1 U281 ( .A1(n835), .A2(n19), .B1(N873), .B2(n256), .ZN(n553) );
  OAI22_X1 U282 ( .A1(n843), .A2(n21), .B1(N881), .B2(n216), .ZN(n577) );
  OAI22_X1 U283 ( .A1(n843), .A2(n21), .B1(N881), .B2(n248), .ZN(n545) );
  OAI22_X1 U284 ( .A1(n833), .A2(n22), .B1(N871), .B2(n226), .ZN(n587) );
  OAI22_X1 U285 ( .A1(n833), .A2(n19), .B1(N871), .B2(n258), .ZN(n555) );
  OAI22_X1 U286 ( .A1(n841), .A2(n21), .B1(N879), .B2(n218), .ZN(n579) );
  OAI22_X1 U287 ( .A1(n841), .A2(n22), .B1(N879), .B2(n250), .ZN(n547) );
  OAI22_X1 U288 ( .A1(n840), .A2(n21), .B1(N878), .B2(n219), .ZN(n580) );
  OAI22_X1 U289 ( .A1(n840), .A2(n24), .B1(N878), .B2(n251), .ZN(n548) );
  OAI22_X1 U290 ( .A1(n848), .A2(n19), .B1(N886), .B2(n211), .ZN(n572) );
  OAI22_X1 U291 ( .A1(n848), .A2(n20), .B1(N886), .B2(n243), .ZN(n540) );
  OAI22_X1 U292 ( .A1(n838), .A2(n21), .B1(N876), .B2(n221), .ZN(n582) );
  OAI22_X1 U293 ( .A1(n838), .A2(n19), .B1(N876), .B2(n253), .ZN(n550) );
  OAI22_X1 U294 ( .A1(n846), .A2(n20), .B1(N884), .B2(n213), .ZN(n574) );
  OAI22_X1 U295 ( .A1(n846), .A2(n24), .B1(N884), .B2(n245), .ZN(n542) );
  OAI22_X1 U296 ( .A1(n836), .A2(n21), .B1(N874), .B2(n223), .ZN(n584) );
  OAI22_X1 U297 ( .A1(n836), .A2(n19), .B1(N874), .B2(n255), .ZN(n552) );
  OAI22_X1 U298 ( .A1(n844), .A2(n21), .B1(N882), .B2(n215), .ZN(n576) );
  OAI22_X1 U299 ( .A1(n844), .A2(n23), .B1(N882), .B2(n247), .ZN(n544) );
  OAI22_X1 U300 ( .A1(n834), .A2(n20), .B1(N872), .B2(n225), .ZN(n586) );
  OAI22_X1 U301 ( .A1(n834), .A2(n19), .B1(N872), .B2(n257), .ZN(n554) );
  OAI22_X1 U302 ( .A1(n842), .A2(n21), .B1(N880), .B2(n217), .ZN(n578) );
  OAI22_X1 U303 ( .A1(n842), .A2(n19), .B1(N880), .B2(n249), .ZN(n546) );
  OAI22_X1 U304 ( .A1(n831), .A2(n22), .B1(N869), .B2(n228), .ZN(n589) );
  OAI22_X1 U305 ( .A1(n831), .A2(n19), .B1(N869), .B2(n260), .ZN(n557) );
  OAI22_X1 U306 ( .A1(n829), .A2(n20), .B1(N867), .B2(n230), .ZN(n591) );
  OAI22_X1 U307 ( .A1(n829), .A2(n20), .B1(N867), .B2(n262), .ZN(n559) );
  OAI22_X1 U308 ( .A1(n827), .A2(n21), .B1(N865), .B2(n232), .ZN(n593) );
  OAI22_X1 U309 ( .A1(n827), .A2(n20), .B1(N865), .B2(n264), .ZN(n561) );
  OAI22_X1 U310 ( .A1(n825), .A2(n21), .B1(N863), .B2(n234), .ZN(n595) );
  OAI22_X1 U311 ( .A1(n825), .A2(n20), .B1(N863), .B2(n266), .ZN(n563) );
  OAI22_X1 U312 ( .A1(n832), .A2(n22), .B1(N870), .B2(n227), .ZN(n588) );
  OAI22_X1 U314 ( .A1(n832), .A2(n19), .B1(N870), .B2(n259), .ZN(n556) );
  OAI22_X1 U315 ( .A1(n830), .A2(n20), .B1(N868), .B2(n229), .ZN(n590) );
  OAI22_X1 U316 ( .A1(n830), .A2(n19), .B1(N868), .B2(n261), .ZN(n558) );
  OAI22_X1 U317 ( .A1(n828), .A2(n24), .B1(N866), .B2(n231), .ZN(n592) );
  OAI22_X1 U318 ( .A1(n828), .A2(n20), .B1(N866), .B2(n263), .ZN(n560) );
  OAI22_X1 U319 ( .A1(n826), .A2(n23), .B1(N864), .B2(n233), .ZN(n594) );
  OAI22_X1 U320 ( .A1(n826), .A2(n20), .B1(N864), .B2(n265), .ZN(n562) );
  INV_X1 U321 ( .A(n428), .ZN(n140) );
  AOI22_X1 U322 ( .A1(gprs_base_addr_o[8]), .A2(n25), .B1(
        warp_pool_wr_data_out[105]), .B2(n39), .ZN(n428) );
  INV_X1 U323 ( .A(n431), .ZN(n157) );
  AOI22_X1 U324 ( .A1(gprs_base_addr_o[5]), .A2(n26), .B1(
        warp_pool_wr_data_out[102]), .B2(n39), .ZN(n431) );
  OAI22_X1 U325 ( .A1(n855), .A2(n20), .B1(N893), .B2(n204), .ZN(n565) );
  OAI22_X1 U326 ( .A1(n855), .A2(n24), .B1(N893), .B2(n236), .ZN(n533) );
  OAI22_X1 U327 ( .A1(n853), .A2(n20), .B1(N891), .B2(n206), .ZN(n567) );
  OAI22_X1 U328 ( .A1(n853), .A2(n21), .B1(N891), .B2(n238), .ZN(n535) );
  OAI22_X1 U329 ( .A1(n851), .A2(n21), .B1(N889), .B2(n208), .ZN(n569) );
  OAI22_X1 U330 ( .A1(n851), .A2(n20), .B1(N889), .B2(n240), .ZN(n537) );
  OAI22_X1 U331 ( .A1(n849), .A2(n21), .B1(N887), .B2(n210), .ZN(n571) );
  OAI22_X1 U332 ( .A1(n849), .A2(n22), .B1(N887), .B2(n242), .ZN(n539) );
  OAI22_X1 U333 ( .A1(n856), .A2(n20), .B1(N894), .B2(n203), .ZN(n564) );
  OAI22_X1 U334 ( .A1(n856), .A2(n19), .B1(N894), .B2(n235), .ZN(n532) );
  OAI22_X1 U335 ( .A1(n854), .A2(n20), .B1(N892), .B2(n205), .ZN(n566) );
  OAI22_X1 U336 ( .A1(n854), .A2(n23), .B1(N892), .B2(n237), .ZN(n534) );
  OAI22_X1 U337 ( .A1(n852), .A2(n21), .B1(N890), .B2(n207), .ZN(n568) );
  OAI22_X1 U338 ( .A1(n852), .A2(n21), .B1(N890), .B2(n239), .ZN(n536) );
  OAI22_X1 U339 ( .A1(n850), .A2(n19), .B1(N888), .B2(n209), .ZN(n570) );
  OAI22_X1 U340 ( .A1(n850), .A2(n20), .B1(N888), .B2(n241), .ZN(n538) );
  OAI22_X1 U341 ( .A1(n486), .A2(n143), .B1(block_num_cnt[1]), .B2(n483), .ZN(
        n811) );
  OAI22_X1 U342 ( .A1(n36), .A2(n40), .B1(n24), .B2(n152), .ZN(n729) );
  OAI22_X1 U343 ( .A1(n37), .A2(n41), .B1(n23), .B2(n153), .ZN(n730) );
  OAI22_X1 U344 ( .A1(n36), .A2(n42), .B1(n22), .B2(n154), .ZN(n731) );
  AND2_X1 U345 ( .A1(warps_per_block_in[0]), .A2(n151), .ZN(n129) );
  OAI22_X1 U346 ( .A1(n202), .A2(n492), .B1(n198), .B2(n510), .ZN(n815) );
  NOR2_X1 U347 ( .A1(n38), .A2(n413), .ZN(n510) );
  OAI22_X1 U348 ( .A1(n37), .A2(n43), .B1(n19), .B2(n155), .ZN(n732) );
  OAI21_X1 U349 ( .B1(n473), .B2(n147), .A(n479), .ZN(n806) );
  OAI21_X1 U350 ( .B1(n473), .B2(n148), .A(n478), .ZN(n805) );
  OAI21_X1 U351 ( .B1(n473), .B2(n149), .A(n477), .ZN(n804) );
  OAI21_X1 U352 ( .B1(n473), .B2(n150), .A(n476), .ZN(n803) );
  OAI21_X1 U353 ( .B1(n473), .B2(n151), .A(n474), .ZN(n802) );
  OAI21_X1 U354 ( .B1(n201), .B2(n492), .A(n493), .ZN(n814) );
  OAI21_X1 U355 ( .B1(n480), .B2(n413), .A(n492), .ZN(n493) );
  OAI21_X1 U356 ( .B1(n831), .B2(n7), .A(n387), .ZN(n699) );
  OAI21_X1 U357 ( .B1(n831), .B2(n10), .A(n386), .ZN(n698) );
  OAI21_X1 U358 ( .B1(n831), .B2(n13), .A(n385), .ZN(n697) );
  OAI21_X1 U359 ( .B1(n831), .B2(n16), .A(n384), .ZN(n696) );
  OAI21_X1 U360 ( .B1(n839), .B2(n8), .A(n355), .ZN(n667) );
  OAI21_X1 U361 ( .B1(n839), .B2(n11), .A(n354), .ZN(n666) );
  OAI21_X1 U362 ( .B1(n839), .B2(n14), .A(n353), .ZN(n665) );
  OAI21_X1 U363 ( .B1(n839), .B2(n17), .A(n352), .ZN(n664) );
  OAI21_X1 U364 ( .B1(n847), .B2(n8), .A(n323), .ZN(n635) );
  OAI21_X1 U365 ( .B1(n847), .B2(n11), .A(n322), .ZN(n634) );
  OAI21_X1 U366 ( .B1(n847), .B2(n14), .A(n321), .ZN(n633) );
  OAI21_X1 U367 ( .B1(n847), .B2(n17), .A(n320), .ZN(n632) );
  OAI21_X1 U368 ( .B1(n829), .B2(n7), .A(n395), .ZN(n707) );
  OAI21_X1 U369 ( .B1(n829), .B2(n10), .A(n394), .ZN(n706) );
  OAI21_X1 U370 ( .B1(n829), .B2(n13), .A(n393), .ZN(n705) );
  OAI21_X1 U371 ( .B1(n829), .B2(n16), .A(n392), .ZN(n704) );
  OAI21_X1 U372 ( .B1(n837), .B2(n8), .A(n363), .ZN(n675) );
  OAI21_X1 U373 ( .B1(n837), .B2(n11), .A(n362), .ZN(n674) );
  OAI21_X1 U374 ( .B1(n837), .B2(n14), .A(n361), .ZN(n673) );
  OAI21_X1 U375 ( .B1(n837), .B2(n17), .A(n360), .ZN(n672) );
  OAI21_X1 U376 ( .B1(n845), .B2(n8), .A(n331), .ZN(n643) );
  OAI21_X1 U377 ( .B1(n845), .B2(n11), .A(n330), .ZN(n642) );
  OAI21_X1 U378 ( .B1(n845), .B2(n14), .A(n329), .ZN(n641) );
  OAI21_X1 U379 ( .B1(n845), .B2(n17), .A(n328), .ZN(n640) );
  OAI21_X1 U380 ( .B1(n827), .B2(n7), .A(n403), .ZN(n715) );
  OAI21_X1 U381 ( .B1(n827), .B2(n10), .A(n402), .ZN(n714) );
  OAI21_X1 U382 ( .B1(n827), .B2(n13), .A(n401), .ZN(n713) );
  OAI21_X1 U383 ( .B1(n827), .B2(n16), .A(n400), .ZN(n712) );
  OAI21_X1 U384 ( .B1(n835), .B2(n7), .A(n371), .ZN(n683) );
  OAI21_X1 U385 ( .B1(n835), .B2(n10), .A(n370), .ZN(n682) );
  OAI21_X1 U386 ( .B1(n835), .B2(n13), .A(n369), .ZN(n681) );
  OAI21_X1 U387 ( .B1(n835), .B2(n16), .A(n368), .ZN(n680) );
  OAI21_X1 U388 ( .B1(n843), .B2(n8), .A(n339), .ZN(n651) );
  OAI21_X1 U389 ( .B1(n843), .B2(n11), .A(n338), .ZN(n650) );
  OAI21_X1 U390 ( .B1(n843), .B2(n14), .A(n337), .ZN(n649) );
  OAI21_X1 U391 ( .B1(n843), .B2(n17), .A(n336), .ZN(n648) );
  OAI21_X1 U392 ( .B1(n825), .B2(n7), .A(n411), .ZN(n723) );
  OAI21_X1 U393 ( .B1(n825), .B2(n10), .A(n410), .ZN(n722) );
  OAI21_X1 U394 ( .B1(n825), .B2(n13), .A(n409), .ZN(n721) );
  OAI21_X1 U395 ( .B1(n825), .B2(n16), .A(n408), .ZN(n720) );
  OAI21_X1 U396 ( .B1(n833), .B2(n7), .A(n379), .ZN(n691) );
  OAI21_X1 U397 ( .B1(n833), .B2(n10), .A(n378), .ZN(n690) );
  OAI21_X1 U398 ( .B1(n833), .B2(n13), .A(n377), .ZN(n689) );
  OAI21_X1 U399 ( .B1(n833), .B2(n16), .A(n376), .ZN(n688) );
  OAI21_X1 U400 ( .B1(n841), .B2(n8), .A(n347), .ZN(n659) );
  OAI21_X1 U401 ( .B1(n841), .B2(n11), .A(n346), .ZN(n658) );
  OAI21_X1 U402 ( .B1(n841), .B2(n14), .A(n345), .ZN(n657) );
  OAI21_X1 U403 ( .B1(n841), .B2(n17), .A(n344), .ZN(n656) );
  OAI21_X1 U404 ( .B1(n832), .B2(n7), .A(n383), .ZN(n695) );
  OAI21_X1 U405 ( .B1(n832), .B2(n10), .A(n382), .ZN(n694) );
  OAI21_X1 U406 ( .B1(n832), .B2(n13), .A(n381), .ZN(n693) );
  OAI21_X1 U407 ( .B1(n832), .B2(n16), .A(n380), .ZN(n692) );
  OAI21_X1 U408 ( .B1(n840), .B2(n8), .A(n351), .ZN(n663) );
  OAI21_X1 U409 ( .B1(n840), .B2(n11), .A(n350), .ZN(n662) );
  OAI21_X1 U410 ( .B1(n840), .B2(n14), .A(n349), .ZN(n661) );
  OAI21_X1 U411 ( .B1(n840), .B2(n17), .A(n348), .ZN(n660) );
  OAI21_X1 U412 ( .B1(n848), .B2(n8), .A(n319), .ZN(n631) );
  OAI21_X1 U413 ( .B1(n848), .B2(n11), .A(n318), .ZN(n630) );
  OAI21_X1 U414 ( .B1(n848), .B2(n14), .A(n317), .ZN(n629) );
  OAI21_X1 U415 ( .B1(n848), .B2(n17), .A(n316), .ZN(n628) );
  OAI21_X1 U416 ( .B1(n830), .B2(n7), .A(n391), .ZN(n703) );
  OAI21_X1 U417 ( .B1(n830), .B2(n10), .A(n390), .ZN(n702) );
  OAI21_X1 U418 ( .B1(n830), .B2(n13), .A(n389), .ZN(n701) );
  OAI21_X1 U419 ( .B1(n830), .B2(n16), .A(n388), .ZN(n700) );
  OAI21_X1 U420 ( .B1(n838), .B2(n8), .A(n359), .ZN(n671) );
  OAI21_X1 U421 ( .B1(n838), .B2(n11), .A(n358), .ZN(n670) );
  OAI21_X1 U422 ( .B1(n838), .B2(n14), .A(n357), .ZN(n669) );
  OAI21_X1 U423 ( .B1(n838), .B2(n17), .A(n356), .ZN(n668) );
  OAI21_X1 U424 ( .B1(n846), .B2(n8), .A(n327), .ZN(n639) );
  OAI21_X1 U425 ( .B1(n846), .B2(n11), .A(n326), .ZN(n638) );
  OAI21_X1 U426 ( .B1(n846), .B2(n14), .A(n325), .ZN(n637) );
  OAI21_X1 U427 ( .B1(n846), .B2(n17), .A(n324), .ZN(n636) );
  OAI21_X1 U428 ( .B1(n828), .B2(n7), .A(n399), .ZN(n711) );
  OAI21_X1 U430 ( .B1(n828), .B2(n10), .A(n398), .ZN(n710) );
  OAI21_X1 U431 ( .B1(n828), .B2(n13), .A(n397), .ZN(n709) );
  OAI21_X1 U432 ( .B1(n828), .B2(n16), .A(n396), .ZN(n708) );
  OAI21_X1 U433 ( .B1(n836), .B2(n7), .A(n367), .ZN(n679) );
  OAI21_X1 U434 ( .B1(n836), .B2(n10), .A(n366), .ZN(n678) );
  OAI21_X1 U435 ( .B1(n836), .B2(n13), .A(n365), .ZN(n677) );
  OAI21_X1 U436 ( .B1(n836), .B2(n16), .A(n364), .ZN(n676) );
  OAI21_X1 U437 ( .B1(n844), .B2(n8), .A(n335), .ZN(n647) );
  OAI21_X1 U438 ( .B1(n844), .B2(n11), .A(n334), .ZN(n646) );
  OAI21_X1 U439 ( .B1(n844), .B2(n14), .A(n333), .ZN(n645) );
  OAI21_X1 U440 ( .B1(n844), .B2(n17), .A(n332), .ZN(n644) );
  OAI21_X1 U441 ( .B1(n826), .B2(n7), .A(n407), .ZN(n719) );
  OAI21_X1 U442 ( .B1(n826), .B2(n10), .A(n406), .ZN(n718) );
  OAI21_X1 U443 ( .B1(n826), .B2(n13), .A(n405), .ZN(n717) );
  OAI21_X1 U444 ( .B1(n826), .B2(n16), .A(n404), .ZN(n716) );
  OAI21_X1 U445 ( .B1(n834), .B2(n7), .A(n375), .ZN(n687) );
  OAI21_X1 U446 ( .B1(n834), .B2(n10), .A(n374), .ZN(n686) );
  OAI21_X1 U447 ( .B1(n834), .B2(n13), .A(n373), .ZN(n685) );
  OAI21_X1 U448 ( .B1(n834), .B2(n16), .A(n372), .ZN(n684) );
  OAI21_X1 U449 ( .B1(n842), .B2(n8), .A(n343), .ZN(n655) );
  OAI21_X1 U450 ( .B1(n842), .B2(n11), .A(n342), .ZN(n654) );
  OAI21_X1 U451 ( .B1(n842), .B2(n14), .A(n341), .ZN(n653) );
  OAI21_X1 U452 ( .B1(n842), .B2(n17), .A(n340), .ZN(n652) );
  OAI21_X1 U453 ( .B1(n38), .B2(n90), .A(n23), .ZN(n771) );
  OAI21_X1 U454 ( .B1(n37), .B2(n78), .A(n23), .ZN(n759) );
  OAI21_X1 U455 ( .B1(n37), .B2(n75), .A(n23), .ZN(n756) );
  OAI21_X1 U456 ( .B1(n37), .B2(n74), .A(n23), .ZN(n755) );
  OAI21_X1 U457 ( .B1(n37), .B2(n73), .A(n23), .ZN(n754) );
  OAI21_X1 U458 ( .B1(n37), .B2(n72), .A(n23), .ZN(n753) );
  OAI21_X1 U459 ( .B1(n36), .B2(n71), .A(n23), .ZN(n752) );
  OAI21_X1 U460 ( .B1(n36), .B2(n70), .A(n23), .ZN(n751) );
  OAI21_X1 U461 ( .B1(n36), .B2(n69), .A(n23), .ZN(n750) );
  OAI21_X1 U462 ( .B1(n36), .B2(n67), .A(n23), .ZN(n748) );
  OAI21_X1 U463 ( .B1(n36), .B2(n115), .A(n20), .ZN(n796) );
  OAI21_X1 U464 ( .B1(n37), .B2(n57), .A(n22), .ZN(n738) );
  OAI21_X1 U465 ( .B1(n36), .B2(n56), .A(n22), .ZN(n737) );
  OAI21_X1 U466 ( .B1(n37), .B2(n55), .A(n20), .ZN(n736) );
  OAI21_X1 U467 ( .B1(n36), .B2(n54), .A(n23), .ZN(n735) );
  OAI21_X1 U468 ( .B1(n37), .B2(n53), .A(n24), .ZN(n734) );
  OAI21_X1 U469 ( .B1(n36), .B2(n116), .A(n23), .ZN(n733) );
  NOR2_X1 U470 ( .A1(block_num_cnt[2]), .A2(n515), .ZN(n514) );
  OAI21_X1 U471 ( .B1(n36), .B2(n109), .A(n21), .ZN(n790) );
  OAI21_X1 U472 ( .B1(n37), .B2(n108), .A(n21), .ZN(n789) );
  OAI21_X1 U473 ( .B1(n36), .B2(n107), .A(n22), .ZN(n788) );
  OAI21_X1 U474 ( .B1(n37), .B2(n106), .A(n24), .ZN(n787) );
  OAI21_X1 U475 ( .B1(n36), .B2(n105), .A(n23), .ZN(n786) );
  OAI21_X1 U476 ( .B1(n37), .B2(n104), .A(n19), .ZN(n785) );
  OAI21_X1 U477 ( .B1(n36), .B2(n103), .A(n19), .ZN(n784) );
  OAI21_X1 U478 ( .B1(n38), .B2(n102), .A(n21), .ZN(n783) );
  OAI21_X1 U479 ( .B1(n38), .B2(n101), .A(n24), .ZN(n782) );
  OAI21_X1 U480 ( .B1(n38), .B2(n100), .A(n23), .ZN(n781) );
  OAI21_X1 U481 ( .B1(n38), .B2(n99), .A(n19), .ZN(n780) );
  OAI21_X1 U482 ( .B1(n38), .B2(n98), .A(n19), .ZN(n779) );
  OAI21_X1 U483 ( .B1(n38), .B2(n97), .A(n19), .ZN(n778) );
  OAI21_X1 U484 ( .B1(n38), .B2(n96), .A(n19), .ZN(n777) );
  OAI21_X1 U485 ( .B1(n38), .B2(n95), .A(n19), .ZN(n776) );
  OAI21_X1 U486 ( .B1(n38), .B2(n94), .A(n23), .ZN(n775) );
  OAI21_X1 U487 ( .B1(n38), .B2(n93), .A(n23), .ZN(n774) );
  OAI21_X1 U488 ( .B1(n38), .B2(n92), .A(n24), .ZN(n773) );
  OAI21_X1 U489 ( .B1(n38), .B2(n91), .A(n23), .ZN(n772) );
  OAI21_X1 U490 ( .B1(n38), .B2(n89), .A(n24), .ZN(n770) );
  OAI21_X1 U491 ( .B1(n38), .B2(n88), .A(n24), .ZN(n769) );
  OAI21_X1 U492 ( .B1(n38), .B2(n87), .A(n24), .ZN(n768) );
  OAI21_X1 U493 ( .B1(n38), .B2(n86), .A(n24), .ZN(n767) );
  OAI21_X1 U494 ( .B1(n38), .B2(n85), .A(n24), .ZN(n766) );
  OAI21_X1 U495 ( .B1(n38), .B2(n84), .A(n24), .ZN(n765) );
  OAI21_X1 U496 ( .B1(n37), .B2(n83), .A(n21), .ZN(n764) );
  OAI21_X1 U497 ( .B1(n37), .B2(n82), .A(n24), .ZN(n763) );
  OAI21_X1 U498 ( .B1(n37), .B2(n81), .A(n24), .ZN(n762) );
  OAI21_X1 U499 ( .B1(n37), .B2(n80), .A(n24), .ZN(n761) );
  OAI21_X1 U500 ( .B1(n37), .B2(n79), .A(n24), .ZN(n760) );
  OAI21_X1 U501 ( .B1(n37), .B2(n77), .A(n24), .ZN(n758) );
  OAI21_X1 U502 ( .B1(n37), .B2(n76), .A(n22), .ZN(n757) );
  OAI21_X1 U503 ( .B1(n36), .B2(n68), .A(n22), .ZN(n749) );
  OAI21_X1 U504 ( .B1(n36), .B2(n66), .A(n22), .ZN(n747) );
  OAI21_X1 U505 ( .B1(n36), .B2(n65), .A(n22), .ZN(n746) );
  OAI21_X1 U506 ( .B1(n37), .B2(n64), .A(n22), .ZN(n745) );
  OAI21_X1 U507 ( .B1(n36), .B2(n63), .A(n22), .ZN(n744) );
  OAI21_X1 U508 ( .B1(n36), .B2(n62), .A(n22), .ZN(n743) );
  OAI21_X1 U509 ( .B1(n36), .B2(n61), .A(n22), .ZN(n742) );
  OAI21_X1 U510 ( .B1(n36), .B2(n60), .A(n22), .ZN(n741) );
  OAI21_X1 U511 ( .B1(n36), .B2(n59), .A(n22), .ZN(n740) );
  OAI21_X1 U512 ( .B1(n36), .B2(n58), .A(n20), .ZN(n739) );
  OAI21_X1 U513 ( .B1(n855), .B2(n9), .A(n291), .ZN(n603) );
  OAI21_X1 U514 ( .B1(n855), .B2(n12), .A(n290), .ZN(n602) );
  OAI21_X1 U515 ( .B1(n855), .B2(n15), .A(n289), .ZN(n601) );
  OAI21_X1 U516 ( .B1(n855), .B2(n18), .A(n288), .ZN(n600) );
  OAI21_X1 U517 ( .B1(n853), .B2(n9), .A(n299), .ZN(n611) );
  OAI21_X1 U518 ( .B1(n853), .B2(n12), .A(n298), .ZN(n610) );
  OAI21_X1 U519 ( .B1(n853), .B2(n15), .A(n297), .ZN(n609) );
  OAI21_X1 U520 ( .B1(n853), .B2(n18), .A(n296), .ZN(n608) );
  OAI21_X1 U521 ( .B1(n851), .B2(n9), .A(n307), .ZN(n619) );
  OAI21_X1 U522 ( .B1(n851), .B2(n12), .A(n306), .ZN(n618) );
  OAI21_X1 U523 ( .B1(n851), .B2(n15), .A(n305), .ZN(n617) );
  OAI21_X1 U524 ( .B1(n851), .B2(n18), .A(n304), .ZN(n616) );
  OAI21_X1 U525 ( .B1(n849), .B2(n9), .A(n315), .ZN(n627) );
  OAI21_X1 U526 ( .B1(n849), .B2(n12), .A(n314), .ZN(n626) );
  OAI21_X1 U527 ( .B1(n849), .B2(n15), .A(n313), .ZN(n625) );
  OAI21_X1 U528 ( .B1(n849), .B2(n18), .A(n312), .ZN(n624) );
  OAI21_X1 U529 ( .B1(n856), .B2(n9), .A(n287), .ZN(n599) );
  OAI21_X1 U530 ( .B1(n856), .B2(n12), .A(n285), .ZN(n598) );
  OAI21_X1 U531 ( .B1(n856), .B2(n15), .A(n283), .ZN(n597) );
  OAI21_X1 U532 ( .B1(n856), .B2(n18), .A(n281), .ZN(n596) );
  OAI21_X1 U533 ( .B1(n854), .B2(n9), .A(n295), .ZN(n607) );
  OAI21_X1 U534 ( .B1(n854), .B2(n12), .A(n294), .ZN(n606) );
  OAI21_X1 U535 ( .B1(n854), .B2(n15), .A(n293), .ZN(n605) );
  OAI21_X1 U536 ( .B1(n854), .B2(n18), .A(n292), .ZN(n604) );
  OAI21_X1 U537 ( .B1(n852), .B2(n9), .A(n303), .ZN(n615) );
  OAI21_X1 U538 ( .B1(n852), .B2(n12), .A(n302), .ZN(n614) );
  OAI21_X1 U539 ( .B1(n852), .B2(n15), .A(n301), .ZN(n613) );
  OAI21_X1 U540 ( .B1(n852), .B2(n18), .A(n300), .ZN(n612) );
  OAI21_X1 U541 ( .B1(n850), .B2(n9), .A(n311), .ZN(n623) );
  OAI21_X1 U542 ( .B1(n850), .B2(n12), .A(n310), .ZN(n622) );
  OAI21_X1 U543 ( .B1(n850), .B2(n15), .A(n309), .ZN(n621) );
  OAI21_X1 U544 ( .B1(n850), .B2(n18), .A(n308), .ZN(n620) );
  OAI21_X1 U545 ( .B1(n145), .B2(n275), .A(n487), .ZN(n810) );
  OAI21_X1 U546 ( .B1(n481), .B2(n141), .A(n482), .ZN(n808) );
  NOR2_X1 U547 ( .A1(n872), .A2(n484), .ZN(n481) );
  OR3_X1 U548 ( .A1(n142), .A2(n143), .A3(n483), .ZN(n482) );
  INV_X1 U549 ( .A(warps_per_block_in[3]), .ZN(n136) );
  INV_X1 U550 ( .A(n494), .ZN(n824) );
  AOI22_X1 U551 ( .A1(N102), .A2(n495), .B1(warps_per_block_cnt[10]), .B2(n496), .ZN(n494) );
  INV_X1 U552 ( .A(n497), .ZN(n823) );
  AOI22_X1 U553 ( .A1(N101), .A2(n495), .B1(warps_per_block_cnt[9]), .B2(n496), 
        .ZN(n497) );
  INV_X1 U554 ( .A(n498), .ZN(n822) );
  AOI22_X1 U555 ( .A1(N100), .A2(n495), .B1(warps_per_block_cnt[8]), .B2(n496), 
        .ZN(n498) );
  INV_X1 U556 ( .A(n499), .ZN(n821) );
  AOI22_X1 U557 ( .A1(N99), .A2(n495), .B1(warps_per_block_cnt[7]), .B2(n496), 
        .ZN(n499) );
  INV_X1 U558 ( .A(n500), .ZN(n820) );
  AOI22_X1 U559 ( .A1(N98), .A2(n495), .B1(warps_per_block_cnt[6]), .B2(n496), 
        .ZN(n500) );
  INV_X1 U560 ( .A(n501), .ZN(n819) );
  AOI22_X1 U561 ( .A1(N97), .A2(n495), .B1(warps_per_block_cnt[5]), .B2(n496), 
        .ZN(n501) );
  INV_X1 U562 ( .A(n507), .ZN(n277) );
  AOI22_X1 U563 ( .A1(N103), .A2(n495), .B1(warps_per_block_cnt[11]), .B2(n496), .ZN(n507) );
  OAI22_X1 U564 ( .A1(n472), .A2(n453), .B1(n273), .B2(n156), .ZN(n798) );
  INV_X1 U565 ( .A(n472), .ZN(n273) );
  NOR2_X1 U566 ( .A1(n274), .A2(n413), .ZN(n472) );
  INV_X1 U567 ( .A(n437), .ZN(n196) );
  AOI22_X1 U568 ( .A1(N78), .A2(n438), .B1(shmem_addr_i[0]), .B2(n439), .ZN(
        n437) );
  INV_X1 U569 ( .A(n440), .ZN(n195) );
  AOI22_X1 U570 ( .A1(N79), .A2(n438), .B1(shmem_addr_i[1]), .B2(n439), .ZN(
        n440) );
  INV_X1 U571 ( .A(n441), .ZN(n194) );
  AOI22_X1 U572 ( .A1(N80), .A2(n438), .B1(shmem_addr_i[2]), .B2(n439), .ZN(
        n441) );
  INV_X1 U573 ( .A(n442), .ZN(n193) );
  AOI22_X1 U574 ( .A1(N81), .A2(n438), .B1(shmem_addr_i[3]), .B2(n439), .ZN(
        n442) );
  INV_X1 U575 ( .A(n443), .ZN(n192) );
  AOI22_X1 U576 ( .A1(N82), .A2(n438), .B1(shmem_addr_i[4]), .B2(n439), .ZN(
        n443) );
  INV_X1 U577 ( .A(n444), .ZN(n191) );
  AOI22_X1 U578 ( .A1(N83), .A2(n438), .B1(shmem_addr_i[5]), .B2(n439), .ZN(
        n444) );
  INV_X1 U579 ( .A(n445), .ZN(n190) );
  AOI22_X1 U580 ( .A1(N84), .A2(n438), .B1(shmem_addr_i[6]), .B2(n439), .ZN(
        n445) );
  INV_X1 U581 ( .A(n446), .ZN(n189) );
  AOI22_X1 U582 ( .A1(N85), .A2(n438), .B1(shmem_addr_i[7]), .B2(n439), .ZN(
        n446) );
  INV_X1 U583 ( .A(n447), .ZN(n188) );
  AOI22_X1 U584 ( .A1(N86), .A2(n438), .B1(shmem_addr_i[8]), .B2(n439), .ZN(
        n447) );
  INV_X1 U585 ( .A(n448), .ZN(n187) );
  AOI22_X1 U586 ( .A1(N87), .A2(n438), .B1(shmem_addr_i[9]), .B2(n439), .ZN(
        n448) );
  INV_X1 U587 ( .A(n449), .ZN(n186) );
  AOI22_X1 U588 ( .A1(N88), .A2(n438), .B1(shmem_addr_i[10]), .B2(n439), .ZN(
        n449) );
  INV_X1 U589 ( .A(n450), .ZN(n185) );
  AOI22_X1 U590 ( .A1(N89), .A2(n438), .B1(shmem_addr_i[11]), .B2(n439), .ZN(
        n450) );
  INV_X1 U591 ( .A(n451), .ZN(n184) );
  AOI22_X1 U592 ( .A1(N90), .A2(n438), .B1(shmem_addr_i[12]), .B2(n439), .ZN(
        n451) );
  INV_X1 U593 ( .A(n509), .ZN(n197) );
  AOI22_X1 U594 ( .A1(warp_generator_state_machine[2]), .A2(n198), .B1(n872), 
        .B2(n508), .ZN(n509) );
  INV_X1 U595 ( .A(n429), .ZN(n144) );
  AOI22_X1 U596 ( .A1(gprs_base_addr_o[7]), .A2(n25), .B1(
        warp_pool_wr_data_out[104]), .B2(n39), .ZN(n429) );
  INV_X1 U729 ( .A(n430), .ZN(n146) );
  AOI22_X1 U730 ( .A1(gprs_base_addr_o[6]), .A2(n25), .B1(
        warp_pool_wr_data_out[103]), .B2(n44), .ZN(n430) );
  INV_X1 U760 ( .A(n432), .ZN(n158) );
  AOI22_X1 U761 ( .A1(gprs_base_addr_o[4]), .A2(n26), .B1(
        warp_pool_wr_data_out[101]), .B2(n45), .ZN(n432) );
  INV_X1 U763 ( .A(n433), .ZN(n159) );
  AOI22_X1 U764 ( .A1(gprs_base_addr_o[3]), .A2(n25), .B1(
        warp_pool_wr_data_out[100]), .B2(n44), .ZN(n433) );
  INV_X1 U765 ( .A(n434), .ZN(n160) );
  AOI22_X1 U766 ( .A1(gprs_base_addr_o[2]), .A2(n26), .B1(
        warp_pool_wr_data_out[99]), .B2(n44), .ZN(n434) );
  OAI22_X1 U767 ( .A1(n412), .A2(n180), .B1(n199), .B2(n271), .ZN(n724) );
  INV_X1 U768 ( .A(warp_id_o[0]), .ZN(n180) );
  INV_X1 U769 ( .A(n436), .ZN(n178) );
  AOI22_X1 U770 ( .A1(gprs_base_addr_o[0]), .A2(n27), .B1(
        warp_pool_wr_data_out[97]), .B2(n44), .ZN(n436) );
  INV_X1 U771 ( .A(n435), .ZN(n161) );
  AOI22_X1 U772 ( .A1(gprs_base_addr_o[1]), .A2(n26), .B1(
        warp_pool_wr_data_out[98]), .B2(n39), .ZN(n435) );
  OAI21_X1 U773 ( .B1(n37), .B2(n114), .A(n22), .ZN(n795) );
  OAI21_X1 U774 ( .B1(n36), .B2(n113), .A(n20), .ZN(n794) );
  OAI21_X1 U775 ( .B1(n37), .B2(n112), .A(n24), .ZN(n793) );
  OAI21_X1 U776 ( .B1(n38), .B2(n111), .A(n23), .ZN(n792) );
  OAI21_X1 U777 ( .B1(n37), .B2(n110), .A(n20), .ZN(n791) );
  INV_X1 U778 ( .A(n459), .ZN(n179) );
  AOI22_X1 U779 ( .A1(n180), .A2(n272), .B1(num_warps_out[0]), .B2(n455), .ZN(
        n459) );
  INV_X1 U780 ( .A(n471), .ZN(n181) );
  AOI22_X1 U781 ( .A1(n51), .A2(warp_pool_addr_out[0]), .B1(n33), .B2(
        warp_id_o[0]), .ZN(n471) );
  INV_X1 U782 ( .A(n466), .ZN(n182) );
  AOI22_X1 U783 ( .A1(n49), .A2(warp_state_addr_out[0]), .B1(n31), .B2(
        warp_id_o[0]), .ZN(n466) );
  INV_X1 U784 ( .A(n427), .ZN(n871) );
  AOI22_X1 U785 ( .A1(n48), .A2(warp_pool_wr_data_out[110]), .B1(n29), .B2(
        shmem_addr_i[0]), .ZN(n427) );
  INV_X1 U786 ( .A(n426), .ZN(n870) );
  AOI22_X1 U787 ( .A1(n47), .A2(warp_pool_wr_data_out[111]), .B1(n29), .B2(
        shmem_addr_i[1]), .ZN(n426) );
  INV_X1 U788 ( .A(n425), .ZN(n869) );
  AOI22_X1 U789 ( .A1(n47), .A2(warp_pool_wr_data_out[112]), .B1(n30), .B2(
        shmem_addr_i[2]), .ZN(n425) );
  INV_X1 U790 ( .A(n424), .ZN(n868) );
  AOI22_X1 U791 ( .A1(n48), .A2(warp_pool_wr_data_out[113]), .B1(n29), .B2(
        shmem_addr_i[3]), .ZN(n424) );
  INV_X1 U792 ( .A(n423), .ZN(n867) );
  AOI22_X1 U793 ( .A1(n46), .A2(warp_pool_wr_data_out[114]), .B1(n28), .B2(
        shmem_addr_i[4]), .ZN(n423) );
  INV_X1 U794 ( .A(n422), .ZN(n866) );
  AOI22_X1 U795 ( .A1(n46), .A2(warp_pool_wr_data_out[115]), .B1(n30), .B2(
        shmem_addr_i[5]), .ZN(n422) );
  INV_X1 U796 ( .A(n421), .ZN(n865) );
  AOI22_X1 U797 ( .A1(n46), .A2(warp_pool_wr_data_out[116]), .B1(n28), .B2(
        shmem_addr_i[6]), .ZN(n421) );
  INV_X1 U798 ( .A(n420), .ZN(n864) );
  AOI22_X1 U799 ( .A1(n47), .A2(warp_pool_wr_data_out[117]), .B1(n30), .B2(
        shmem_addr_i[7]), .ZN(n420) );
  INV_X1 U800 ( .A(n419), .ZN(n863) );
  AOI22_X1 U801 ( .A1(n45), .A2(warp_pool_wr_data_out[118]), .B1(n28), .B2(
        shmem_addr_i[8]), .ZN(n419) );
  INV_X1 U802 ( .A(n418), .ZN(n862) );
  AOI22_X1 U803 ( .A1(n47), .A2(warp_pool_wr_data_out[119]), .B1(n28), .B2(
        shmem_addr_i[9]), .ZN(n418) );
  INV_X1 U804 ( .A(n417), .ZN(n861) );
  AOI22_X1 U805 ( .A1(n45), .A2(warp_pool_wr_data_out[120]), .B1(n27), .B2(
        shmem_addr_i[10]), .ZN(n417) );
  INV_X1 U806 ( .A(n416), .ZN(n860) );
  AOI22_X1 U807 ( .A1(n46), .A2(warp_pool_wr_data_out[121]), .B1(n29), .B2(
        shmem_addr_i[11]), .ZN(n416) );
  INV_X1 U808 ( .A(n415), .ZN(n859) );
  AOI22_X1 U809 ( .A1(n45), .A2(warp_pool_wr_data_out[122]), .B1(n27), .B2(
        shmem_addr_i[12]), .ZN(n415) );
  INV_X1 U810 ( .A(n414), .ZN(n858) );
  AOI22_X1 U811 ( .A1(n48), .A2(warp_pool_wr_data_out[123]), .B1(n27), .B2(
        shmem_addr_i[13]), .ZN(n414) );
  INV_X1 U812 ( .A(n34), .ZN(n23) );
  INV_X1 U813 ( .A(n119), .ZN(n122) );
  INV_X1 U814 ( .A(n119), .ZN(n123) );
  INV_X1 U815 ( .A(n119), .ZN(n124) );
  INV_X1 U816 ( .A(n119), .ZN(n125) );
  INV_X1 U817 ( .A(n120), .ZN(n126) );
  INV_X1 U818 ( .A(n120), .ZN(n127) );
  XOR2_X1 U819 ( .A(\add_155/carry[4] ), .B(warp_id_o[4]), .Z(N257) );
  OR4_X1 U820 ( .A1(warps_per_block_cnt[7]), .A2(warps_per_block_cnt[6]), .A3(
        warps_per_block_cnt[9]), .A4(warps_per_block_cnt[8]), .ZN(n135) );
  AND2_X1 U821 ( .A1(n150), .A2(n129), .ZN(n128) );
  OAI222_X1 U822 ( .A1(n129), .A2(n150), .B1(warps_per_block_in[1]), .B2(n128), 
        .C1(warps_per_block_in[2]), .C2(n149), .ZN(n130) );
  AOI221_X1 U823 ( .B1(n149), .B2(warps_per_block_in[2]), .C1(n148), .C2(
        warps_per_block_in[3]), .A(n138), .ZN(n131) );
  AOI221_X1 U824 ( .B1(n136), .B2(warps_per_block_cnt[3]), .C1(n137), .C2(
        warps_per_block_cnt[4]), .A(n131), .ZN(n132) );
  AOI221_X1 U825 ( .B1(n147), .B2(warps_per_block_in[4]), .C1(n2), .C2(
        warps_per_block_in[5]), .A(n132), .ZN(n133) );
  OAI21_X1 U826 ( .B1(warps_per_block_in[5]), .B2(n2), .A(n139), .ZN(n134) );
  NOR4_X1 U827 ( .A1(n135), .A2(n134), .A3(warps_per_block_cnt[11]), .A4(
        warps_per_block_cnt[10]), .ZN(N62) );
  NAND2_X1 U828 ( .A1(n413), .A2(n126), .ZN(n412) );
endmodule





module warp_id_calc_1_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [8:0] A;
  input [8:0] B;
  output [17:0] PRODUCT;
  input TC;
  wire   \ab[8><0] , \ab[7><1] , \ab[7><0] , \ab[6><2] , \ab[6><1] ,
         \ab[6><0] , \ab[5><3] , \ab[5><2] , \ab[5><1] , \ab[5><0] ,
         \ab[4><4] , \ab[4><3] , \ab[4><2] , \ab[4><1] , \ab[4><0] ,
         \ab[3><5] , \ab[3><4] , \ab[3><3] , \ab[3><2] , \ab[3><1] ,
         \ab[3><0] , \ab[2><6] , \ab[2><5] , \ab[2><4] , \ab[2><3] ,
         \ab[2><2] , \ab[2><1] , \ab[2><0] , \ab[1><7] , \ab[1><6] ,
         \ab[1><5] , \ab[1><4] , \ab[1><3] , \ab[1><2] , \ab[1><1] ,
         \ab[1><0] , \ab[0><8] , \ab[0><7] , \ab[0><6] , \ab[0><5] ,
         \ab[0><4] , \ab[0><3] , \ab[0><2] , \ab[0><1] , \CARRYB[7><0] ,
         \CARRYB[6><1] , \CARRYB[6><0] , \CARRYB[5><2] , \CARRYB[5><1] ,
         \CARRYB[5><0] , \CARRYB[4><3] , \CARRYB[4><2] , \CARRYB[4><1] ,
         \CARRYB[4><0] , \CARRYB[3><4] , \CARRYB[3><3] , \CARRYB[3><2] ,
         \CARRYB[3><1] , \CARRYB[3><0] , \CARRYB[2><5] , \CARRYB[2><4] ,
         \CARRYB[2><3] , \CARRYB[2><2] , \CARRYB[2><1] , \CARRYB[2><0] ,
         \SUMB[7><1] , \SUMB[6><2] , \SUMB[6><1] , \SUMB[5><3] , \SUMB[5><2] ,
         \SUMB[5><1] , \SUMB[4><4] , \SUMB[4><3] , \SUMB[4><2] , \SUMB[4><1] ,
         \SUMB[3><5] , \SUMB[3><4] , \SUMB[3><3] , \SUMB[3><2] , \SUMB[3><1] ,
         \SUMB[2><6] , \SUMB[2><5] , \SUMB[2><4] , \SUMB[2><3] , \SUMB[2><2] ,
         \SUMB[2><1] , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34;

  FA_X1 S4_0 ( .A(\ab[8><0] ), .B(\CARRYB[7><0] ), .CI(\SUMB[7><1] ), .S(
        PRODUCT[8]) );
  FA_X1 S1_7_0 ( .A(\ab[7><0] ), .B(\CARRYB[6><0] ), .CI(\SUMB[6><1] ), .CO(
        \CARRYB[7><0] ), .S(PRODUCT[7]) );
  FA_X1 S2_7_1 ( .A(\ab[7><1] ), .B(\CARRYB[6><1] ), .CI(\SUMB[6><2] ), .S(
        \SUMB[7><1] ) );
  FA_X1 S1_6_0 ( .A(\ab[6><0] ), .B(\CARRYB[5><0] ), .CI(\SUMB[5><1] ), .CO(
        \CARRYB[6><0] ), .S(PRODUCT[6]) );
  FA_X1 S2_6_1 ( .A(\ab[6><1] ), .B(\CARRYB[5><1] ), .CI(\SUMB[5><2] ), .CO(
        \CARRYB[6><1] ), .S(\SUMB[6><1] ) );
  FA_X1 S2_6_2 ( .A(\ab[6><2] ), .B(\CARRYB[5><2] ), .CI(\SUMB[5><3] ), .S(
        \SUMB[6><2] ) );
  FA_X1 S1_5_0 ( .A(\ab[5><0] ), .B(\CARRYB[4><0] ), .CI(\SUMB[4><1] ), .CO(
        \CARRYB[5><0] ), .S(PRODUCT[5]) );
  FA_X1 S2_5_1 ( .A(\ab[5><1] ), .B(\CARRYB[4><1] ), .CI(\SUMB[4><2] ), .CO(
        \CARRYB[5><1] ), .S(\SUMB[5><1] ) );
  FA_X1 S2_5_2 ( .A(\ab[5><2] ), .B(\CARRYB[4><2] ), .CI(\SUMB[4><3] ), .CO(
        \CARRYB[5><2] ), .S(\SUMB[5><2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5><3] ), .B(\CARRYB[4><3] ), .CI(\SUMB[4><4] ), .S(
        \SUMB[5><3] ) );
  FA_X1 S1_4_0 ( .A(\ab[4><0] ), .B(\CARRYB[3><0] ), .CI(\SUMB[3><1] ), .CO(
        \CARRYB[4><0] ), .S(PRODUCT[4]) );
  FA_X1 S2_4_1 ( .A(\ab[4><1] ), .B(\CARRYB[3><1] ), .CI(\SUMB[3><2] ), .CO(
        \CARRYB[4><1] ), .S(\SUMB[4><1] ) );
  FA_X1 S2_4_2 ( .A(\ab[4><2] ), .B(\CARRYB[3><2] ), .CI(\SUMB[3><3] ), .CO(
        \CARRYB[4><2] ), .S(\SUMB[4><2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4><3] ), .B(\CARRYB[3><3] ), .CI(\SUMB[3><4] ), .CO(
        \CARRYB[4><3] ), .S(\SUMB[4><3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4><4] ), .B(\CARRYB[3><4] ), .CI(\SUMB[3><5] ), .S(
        \SUMB[4><4] ) );
  FA_X1 S1_3_0 ( .A(\ab[3><0] ), .B(\CARRYB[2><0] ), .CI(\SUMB[2><1] ), .CO(
        \CARRYB[3><0] ), .S(PRODUCT[3]) );
  FA_X1 S2_3_1 ( .A(\ab[3><1] ), .B(\CARRYB[2><1] ), .CI(\SUMB[2><2] ), .CO(
        \CARRYB[3><1] ), .S(\SUMB[3><1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3><2] ), .B(\CARRYB[2><2] ), .CI(\SUMB[2><3] ), .CO(
        \CARRYB[3><2] ), .S(\SUMB[3><2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3><3] ), .B(\CARRYB[2><3] ), .CI(\SUMB[2><4] ), .CO(
        \CARRYB[3><3] ), .S(\SUMB[3><3] ) );
  FA_X1 S2_3_4 ( .A(\ab[3><4] ), .B(\CARRYB[2><4] ), .CI(\SUMB[2><5] ), .CO(
        \CARRYB[3><4] ), .S(\SUMB[3><4] ) );
  FA_X1 S2_3_5 ( .A(\ab[3><5] ), .B(\CARRYB[2><5] ), .CI(\SUMB[2><6] ), .S(
        \SUMB[3><5] ) );
  FA_X1 S1_2_0 ( .A(\ab[2><0] ), .B(n8), .CI(n14), .CO(\CARRYB[2><0] ), .S(
        PRODUCT[2]) );
  FA_X1 S2_2_1 ( .A(\ab[2><1] ), .B(n7), .CI(n13), .CO(\CARRYB[2><1] ), .S(
        \SUMB[2><1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2><2] ), .B(n6), .CI(n12), .CO(\CARRYB[2><2] ), .S(
        \SUMB[2><2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2><3] ), .B(n5), .CI(n11), .CO(\CARRYB[2><3] ), .S(
        \SUMB[2><3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2><4] ), .B(n4), .CI(n10), .CO(\CARRYB[2><4] ), .S(
        \SUMB[2><4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2><5] ), .B(n3), .CI(n9), .CO(\CARRYB[2><5] ), .S(
        \SUMB[2><5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2><6] ), .B(n2), .CI(n15), .S(\SUMB[2><6] ) );
  AND2_X1 U2 ( .A1(\ab[0><7] ), .A2(\ab[1><6] ), .ZN(n2) );
  AND2_X1 U3 ( .A1(\ab[0><6] ), .A2(\ab[1><5] ), .ZN(n3) );
  AND2_X1 U4 ( .A1(\ab[0><5] ), .A2(\ab[1><4] ), .ZN(n4) );
  AND2_X1 U5 ( .A1(\ab[0><4] ), .A2(\ab[1><3] ), .ZN(n5) );
  AND2_X1 U6 ( .A1(\ab[0><3] ), .A2(\ab[1><2] ), .ZN(n6) );
  AND2_X1 U7 ( .A1(\ab[0><2] ), .A2(\ab[1><1] ), .ZN(n7) );
  AND2_X1 U8 ( .A1(\ab[0><1] ), .A2(\ab[1><0] ), .ZN(n8) );
  XOR2_X1 U9 ( .A(\ab[1><6] ), .B(\ab[0><7] ), .Z(n9) );
  XOR2_X1 U10 ( .A(\ab[1><5] ), .B(\ab[0><6] ), .Z(n10) );
  XOR2_X1 U11 ( .A(\ab[1><4] ), .B(\ab[0><5] ), .Z(n11) );
  XOR2_X1 U12 ( .A(\ab[1><3] ), .B(\ab[0><4] ), .Z(n12) );
  XOR2_X1 U13 ( .A(\ab[1><2] ), .B(\ab[0><3] ), .Z(n13) );
  XOR2_X1 U14 ( .A(\ab[1><1] ), .B(\ab[0><2] ), .Z(n14) );
  XOR2_X1 U15 ( .A(\ab[1><7] ), .B(\ab[0><8] ), .Z(n15) );
  XOR2_X1 U16 ( .A(\ab[1><0] ), .B(\ab[0><1] ), .Z(PRODUCT[1]) );
  INV_X1 U17 ( .A(A[8]), .ZN(n17) );
  INV_X1 U18 ( .A(A[7]), .ZN(n18) );
  INV_X1 U19 ( .A(A[6]), .ZN(n19) );
  INV_X1 U20 ( .A(A[5]), .ZN(n20) );
  INV_X1 U21 ( .A(A[0]), .ZN(n25) );
  INV_X1 U22 ( .A(A[1]), .ZN(n24) );
  INV_X1 U23 ( .A(A[2]), .ZN(n23) );
  INV_X1 U24 ( .A(A[3]), .ZN(n22) );
  INV_X1 U25 ( .A(A[4]), .ZN(n21) );
  INV_X1 U26 ( .A(B[8]), .ZN(n26) );
  INV_X1 U27 ( .A(B[0]), .ZN(n34) );
  INV_X1 U28 ( .A(B[1]), .ZN(n33) );
  INV_X1 U29 ( .A(B[2]), .ZN(n32) );
  INV_X1 U30 ( .A(B[3]), .ZN(n31) );
  INV_X1 U31 ( .A(B[4]), .ZN(n30) );
  INV_X1 U32 ( .A(B[5]), .ZN(n29) );
  INV_X1 U33 ( .A(B[6]), .ZN(n28) );
  INV_X1 U34 ( .A(B[7]), .ZN(n27) );
  NOR2_X1 U35 ( .A1(n17), .A2(n34), .ZN(\ab[8><0] ) );
  NOR2_X1 U36 ( .A1(n33), .A2(n18), .ZN(\ab[7><1] ) );
  NOR2_X1 U37 ( .A1(n34), .A2(n18), .ZN(\ab[7><0] ) );
  NOR2_X1 U38 ( .A1(n32), .A2(n19), .ZN(\ab[6><2] ) );
  NOR2_X1 U39 ( .A1(n33), .A2(n19), .ZN(\ab[6><1] ) );
  NOR2_X1 U40 ( .A1(n34), .A2(n19), .ZN(\ab[6><0] ) );
  NOR2_X1 U41 ( .A1(n31), .A2(n20), .ZN(\ab[5><3] ) );
  NOR2_X1 U42 ( .A1(n32), .A2(n20), .ZN(\ab[5><2] ) );
  NOR2_X1 U43 ( .A1(n33), .A2(n20), .ZN(\ab[5><1] ) );
  NOR2_X1 U44 ( .A1(n34), .A2(n20), .ZN(\ab[5><0] ) );
  NOR2_X1 U45 ( .A1(n30), .A2(n21), .ZN(\ab[4><4] ) );
  NOR2_X1 U46 ( .A1(n31), .A2(n21), .ZN(\ab[4><3] ) );
  NOR2_X1 U47 ( .A1(n32), .A2(n21), .ZN(\ab[4><2] ) );
  NOR2_X1 U48 ( .A1(n33), .A2(n21), .ZN(\ab[4><1] ) );
  NOR2_X1 U49 ( .A1(n34), .A2(n21), .ZN(\ab[4><0] ) );
  NOR2_X1 U50 ( .A1(n29), .A2(n22), .ZN(\ab[3><5] ) );
  NOR2_X1 U51 ( .A1(n30), .A2(n22), .ZN(\ab[3><4] ) );
  NOR2_X1 U52 ( .A1(n31), .A2(n22), .ZN(\ab[3><3] ) );
  NOR2_X1 U53 ( .A1(n32), .A2(n22), .ZN(\ab[3><2] ) );
  NOR2_X1 U54 ( .A1(n33), .A2(n22), .ZN(\ab[3><1] ) );
  NOR2_X1 U55 ( .A1(n34), .A2(n22), .ZN(\ab[3><0] ) );
  NOR2_X1 U56 ( .A1(n28), .A2(n23), .ZN(\ab[2><6] ) );
  NOR2_X1 U57 ( .A1(n29), .A2(n23), .ZN(\ab[2><5] ) );
  NOR2_X1 U58 ( .A1(n30), .A2(n23), .ZN(\ab[2><4] ) );
  NOR2_X1 U59 ( .A1(n31), .A2(n23), .ZN(\ab[2><3] ) );
  NOR2_X1 U60 ( .A1(n32), .A2(n23), .ZN(\ab[2><2] ) );
  NOR2_X1 U61 ( .A1(n33), .A2(n23), .ZN(\ab[2><1] ) );
  NOR2_X1 U62 ( .A1(n34), .A2(n23), .ZN(\ab[2><0] ) );
  NOR2_X1 U63 ( .A1(n27), .A2(n24), .ZN(\ab[1><7] ) );
  NOR2_X1 U64 ( .A1(n28), .A2(n24), .ZN(\ab[1><6] ) );
  NOR2_X1 U65 ( .A1(n29), .A2(n24), .ZN(\ab[1><5] ) );
  NOR2_X1 U66 ( .A1(n30), .A2(n24), .ZN(\ab[1><4] ) );
  NOR2_X1 U67 ( .A1(n31), .A2(n24), .ZN(\ab[1><3] ) );
  NOR2_X1 U68 ( .A1(n32), .A2(n24), .ZN(\ab[1><2] ) );
  NOR2_X1 U69 ( .A1(n33), .A2(n24), .ZN(\ab[1><1] ) );
  NOR2_X1 U70 ( .A1(n34), .A2(n24), .ZN(\ab[1><0] ) );
  NOR2_X1 U71 ( .A1(n26), .A2(n25), .ZN(\ab[0><8] ) );
  NOR2_X1 U72 ( .A1(n27), .A2(n25), .ZN(\ab[0><7] ) );
  NOR2_X1 U73 ( .A1(n28), .A2(n25), .ZN(\ab[0><6] ) );
  NOR2_X1 U74 ( .A1(n29), .A2(n25), .ZN(\ab[0><5] ) );
  NOR2_X1 U75 ( .A1(n30), .A2(n25), .ZN(\ab[0><4] ) );
  NOR2_X1 U76 ( .A1(n31), .A2(n25), .ZN(\ab[0><3] ) );
  NOR2_X1 U77 ( .A1(n32), .A2(n25), .ZN(\ab[0><2] ) );
  NOR2_X1 U78 ( .A1(n33), .A2(n25), .ZN(\ab[0><1] ) );
  NOR2_X1 U79 ( .A1(n34), .A2(n25), .ZN(PRODUCT[0]) );
endmodule


module warp_id_calc_1_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [3:0] A;
  input [5:0] B;
  output [9:0] PRODUCT;
  input TC;
  wire   \ab[3><5] , \ab[3><4] , \ab[3><3] , \ab[3><2] , \ab[3><1] ,
         \ab[3><0] , \ab[2><5] , \ab[2><4] , \ab[2><3] , \ab[2><2] ,
         \ab[2><1] , \ab[2><0] , \ab[1><5] , \ab[1><4] , \ab[1><3] ,
         \ab[1><2] , \ab[1><1] , \ab[1><0] , \ab[0><5] , \ab[0><4] ,
         \ab[0><3] , \ab[0><2] , \ab[0><1] , \CARRYB[3><4] , \CARRYB[3><3] ,
         \CARRYB[3><2] , \CARRYB[3><1] , \CARRYB[3><0] , \CARRYB[2><4] ,
         \CARRYB[2><3] , \CARRYB[2><2] , \CARRYB[2><1] , \CARRYB[2><0] ,
         \SUMB[3><4] , \SUMB[3><3] , \SUMB[3><2] , \SUMB[3><1] , \SUMB[2><4] ,
         \SUMB[2><3] , \SUMB[2><2] , \SUMB[2><1] , n2, n3, n4, n5, n6, n7, n8,
         n9, n11, n12, n14, n15, n16, n17, n18, n19, n20, n21, n22, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50;

  FA_X1 S4_0 ( .A(\ab[3><0] ), .B(\CARRYB[2><0] ), .CI(\SUMB[2><1] ), .CO(
        \CARRYB[3><0] ), .S(PRODUCT[3]) );
  FA_X1 S4_1 ( .A(\ab[3><1] ), .B(\CARRYB[2><1] ), .CI(\SUMB[2><2] ), .CO(
        \CARRYB[3><1] ), .S(\SUMB[3><1] ) );
  FA_X1 S4_2 ( .A(\ab[3><2] ), .B(\CARRYB[2><2] ), .CI(\SUMB[2><3] ), .CO(
        \CARRYB[3><2] ), .S(\SUMB[3><2] ) );
  FA_X1 S4_3 ( .A(\ab[3><3] ), .B(\CARRYB[2><3] ), .CI(\SUMB[2><4] ), .CO(
        \CARRYB[3><3] ), .S(\SUMB[3><3] ) );
  FA_X1 S5_4 ( .A(\ab[3><4] ), .B(\CARRYB[2><4] ), .CI(\ab[2><5] ), .CO(
        \CARRYB[3><4] ), .S(\SUMB[3><4] ) );
  FA_X1 S1_2_0 ( .A(\ab[2><0] ), .B(n12), .CI(n5), .CO(\CARRYB[2><0] ), .S(
        PRODUCT[2]) );
  FA_X1 S2_2_1 ( .A(\ab[2><1] ), .B(n4), .CI(n9), .CO(\CARRYB[2><1] ), .S(
        \SUMB[2><1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2><2] ), .B(n3), .CI(n8), .CO(\CARRYB[2><2] ), .S(
        \SUMB[2><2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2><3] ), .B(n2), .CI(n7), .CO(\CARRYB[2><3] ), .S(
        \SUMB[2><3] ) );
  FA_X1 S3_2_4 ( .A(\ab[2><4] ), .B(n6), .CI(\ab[1><5] ), .CO(\CARRYB[2><4] ), 
        .S(\SUMB[2><4] ) );
  AND2_X1 U2 ( .A1(\ab[0><4] ), .A2(\ab[1><3] ), .ZN(n2) );
  AND2_X1 U3 ( .A1(\ab[0><3] ), .A2(\ab[1><2] ), .ZN(n3) );
  AND2_X1 U4 ( .A1(\ab[0><2] ), .A2(\ab[1><1] ), .ZN(n4) );
  XOR2_X1 U5 ( .A(\ab[1><1] ), .B(\ab[0><2] ), .Z(n5) );
  AND2_X1 U6 ( .A1(\ab[0><5] ), .A2(\ab[1><4] ), .ZN(n6) );
  XOR2_X1 U7 ( .A(\ab[1><4] ), .B(\ab[0><5] ), .Z(n7) );
  XOR2_X1 U8 ( .A(\ab[1><3] ), .B(\ab[0><4] ), .Z(n8) );
  XOR2_X1 U9 ( .A(\ab[1><2] ), .B(\ab[0><3] ), .Z(n9) );
  XOR2_X1 U10 ( .A(\CARRYB[3><0] ), .B(\SUMB[3><1] ), .Z(PRODUCT[4]) );
  OR2_X1 U11 ( .A1(n16), .A2(n14), .ZN(n11) );
  AND2_X1 U12 ( .A1(\ab[0><1] ), .A2(\ab[1><0] ), .ZN(n12) );
  INV_X1 U13 ( .A(n31), .ZN(n39) );
  INV_X1 U14 ( .A(n33), .ZN(n40) );
  INV_X1 U15 ( .A(n24), .ZN(n37) );
  INV_X1 U16 ( .A(n26), .ZN(n38) );
  XNOR2_X1 U17 ( .A(n22), .B(n36), .ZN(PRODUCT[9]) );
  AND2_X1 U18 ( .A1(n24), .A2(n11), .ZN(PRODUCT[5]) );
  XOR2_X1 U19 ( .A(\CARRYB[3><1] ), .B(\SUMB[3><2] ), .Z(n14) );
  XOR2_X1 U20 ( .A(\CARRYB[3><4] ), .B(\ab[3><5] ), .Z(n15) );
  AND2_X1 U21 ( .A1(\CARRYB[3><0] ), .A2(\SUMB[3><1] ), .ZN(n16) );
  AND2_X1 U22 ( .A1(\CARRYB[3><2] ), .A2(\SUMB[3><3] ), .ZN(n17) );
  XOR2_X1 U23 ( .A(\CARRYB[3><3] ), .B(\SUMB[3><4] ), .Z(n18) );
  AND2_X1 U24 ( .A1(\CARRYB[3><1] ), .A2(\SUMB[3><2] ), .ZN(n19) );
  AND2_X1 U25 ( .A1(\CARRYB[3><3] ), .A2(\SUMB[3><4] ), .ZN(n20) );
  XOR2_X1 U26 ( .A(\CARRYB[3><2] ), .B(\SUMB[3><3] ), .Z(n21) );
  AND2_X1 U27 ( .A1(\CARRYB[3><4] ), .A2(\ab[3><5] ), .ZN(n22) );
  INV_X1 U28 ( .A(B[2]), .ZN(n48) );
  INV_X1 U29 ( .A(B[4]), .ZN(n46) );
  INV_X1 U30 ( .A(B[3]), .ZN(n47) );
  INV_X1 U31 ( .A(A[0]), .ZN(n44) );
  INV_X1 U32 ( .A(A[1]), .ZN(n41) );
  INV_X1 U33 ( .A(A[2]), .ZN(n42) );
  INV_X1 U34 ( .A(B[1]), .ZN(n49) );
  INV_X1 U35 ( .A(B[0]), .ZN(n50) );
  XOR2_X1 U36 ( .A(\ab[1><0] ), .B(\ab[0><1] ), .Z(PRODUCT[1]) );
  INV_X1 U37 ( .A(B[5]), .ZN(n45) );
  INV_X1 U38 ( .A(A[3]), .ZN(n43) );
  NAND2_X1 U39 ( .A1(n16), .A2(n14), .ZN(n24) );
  NOR2_X1 U40 ( .A1(n19), .A2(n21), .ZN(n26) );
  AND2_X1 U41 ( .A1(n19), .A2(n21), .ZN(n27) );
  NOR2_X1 U42 ( .A1(n26), .A2(n27), .ZN(n25) );
  XOR2_X1 U43 ( .A(n37), .B(n25), .Z(PRODUCT[6]) );
  NAND2_X1 U44 ( .A1(n17), .A2(n18), .ZN(n29) );
  NOR2_X1 U45 ( .A1(n17), .A2(n18), .ZN(n31) );
  NAND2_X1 U46 ( .A1(n29), .A2(n39), .ZN(n28) );
  AOI21_X1 U47 ( .B1(n38), .B2(n37), .A(n27), .ZN(n30) );
  XOR2_X1 U48 ( .A(n28), .B(n30), .Z(PRODUCT[7]) );
  OAI21_X1 U49 ( .B1(n31), .B2(n30), .A(n29), .ZN(n35) );
  NOR2_X1 U50 ( .A1(n20), .A2(n15), .ZN(n33) );
  AND2_X1 U51 ( .A1(n20), .A2(n15), .ZN(n34) );
  NOR2_X1 U52 ( .A1(n33), .A2(n34), .ZN(n32) );
  XOR2_X1 U53 ( .A(n35), .B(n32), .Z(PRODUCT[8]) );
  AOI21_X1 U54 ( .B1(n35), .B2(n40), .A(n34), .ZN(n36) );
  NOR2_X1 U55 ( .A1(n43), .A2(n45), .ZN(\ab[3><5] ) );
  NOR2_X1 U56 ( .A1(n43), .A2(n46), .ZN(\ab[3><4] ) );
  NOR2_X1 U57 ( .A1(n43), .A2(n47), .ZN(\ab[3><3] ) );
  NOR2_X1 U58 ( .A1(n43), .A2(n48), .ZN(\ab[3><2] ) );
  NOR2_X1 U59 ( .A1(n43), .A2(n49), .ZN(\ab[3><1] ) );
  NOR2_X1 U60 ( .A1(n43), .A2(n50), .ZN(\ab[3><0] ) );
  NOR2_X1 U61 ( .A1(n45), .A2(n42), .ZN(\ab[2><5] ) );
  NOR2_X1 U62 ( .A1(n46), .A2(n42), .ZN(\ab[2><4] ) );
  NOR2_X1 U63 ( .A1(n47), .A2(n42), .ZN(\ab[2><3] ) );
  NOR2_X1 U64 ( .A1(n48), .A2(n42), .ZN(\ab[2><2] ) );
  NOR2_X1 U65 ( .A1(n49), .A2(n42), .ZN(\ab[2><1] ) );
  NOR2_X1 U66 ( .A1(n50), .A2(n42), .ZN(\ab[2><0] ) );
  NOR2_X1 U67 ( .A1(n45), .A2(n41), .ZN(\ab[1><5] ) );
  NOR2_X1 U68 ( .A1(n46), .A2(n41), .ZN(\ab[1><4] ) );
  NOR2_X1 U69 ( .A1(n47), .A2(n41), .ZN(\ab[1><3] ) );
  NOR2_X1 U70 ( .A1(n48), .A2(n41), .ZN(\ab[1><2] ) );
  NOR2_X1 U71 ( .A1(n49), .A2(n41), .ZN(\ab[1><1] ) );
  NOR2_X1 U72 ( .A1(n50), .A2(n41), .ZN(\ab[1><0] ) );
  NOR2_X1 U73 ( .A1(n45), .A2(n44), .ZN(\ab[0><5] ) );
  NOR2_X1 U74 ( .A1(n46), .A2(n44), .ZN(\ab[0><4] ) );
  NOR2_X1 U75 ( .A1(n47), .A2(n44), .ZN(\ab[0><3] ) );
  NOR2_X1 U76 ( .A1(n48), .A2(n44), .ZN(\ab[0><2] ) );
  NOR2_X1 U77 ( .A1(n49), .A2(n44), .ZN(\ab[0><1] ) );
  NOR2_X1 U78 ( .A1(n50), .A2(n44), .ZN(PRODUCT[0]) );
endmodule


module warp_id_calc ( clk, reset, en, block_num_in, gprs_size_in, 
        warp_num_in, warps_per_block_in, data_valid_out, gprs_base_addr_out, 
        warp_id_out );
  input [3:0] block_num_in;
  input [8:0] gprs_size_in;
  input [4:0] warp_num_in;
  input [5:0] warps_per_block_in;
  output [8:0] gprs_base_addr_out;
  output [4:0] warp_id_out;
  input clk, reset, en;
  output data_valid_out;
  wire   N9, N8, N7, N6, N5, N4, N3, N2, N1, N0, \rem_36/u_div/PartRem[4><5] ,
         \rem_36/u_div/PartRem[4><4] , \rem_36/u_div/PartRem[4><3] ,
         \rem_36/u_div/PartRem[4><2] , \rem_36/u_div/PartRem[3><5] ,
         \rem_36/u_div/PartRem[3><4] , \rem_36/u_div/PartRem[3><3] ,
         \rem_36/u_div/PartRem[3><2] , \rem_36/u_div/PartRem[2><5] ,
         \rem_36/u_div/PartRem[2><4] , \rem_36/u_div/PartRem[2><3] ,
         \rem_36/u_div/PartRem[2><2] , \rem_36/u_div/PartRem[1><5] ,
         \rem_36/u_div/PartRem[1><4] , \rem_36/u_div/PartRem[1><3] ,
         \rem_36/u_div/PartRem[1><2] , \add_35/carry[9] , \add_35/carry[8] ,
         \add_35/carry[7] , \add_35/carry[6] , \add_35/carry[5] ,
         \add_35/carry[4] , \add_35/carry[3] , \add_35/carry[2] ,
         \add_35/carry[1] ;
  wire   [9:0] q_res;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8;
  assign data_valid_out = 1'b1;

  warp_id_calc_1_DW02_mult_1 mult_39 ( .A({q_res[8:1], warp_id_out[0]}), .B(
        gprs_size_in), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, gprs_base_addr_out})
         );
  warp_id_calc_1_DW02_mult_0 mult_35 ( .A(block_num_in), .B(warps_per_block_in), .TC(1'b0), .PRODUCT({N9, N8, N7, N6, N5, N4, N3, N2, N1, N0}) );
  FA_X1 \add_35/U1_1  ( .A(N1), .B(warp_num_in[1]), .CI(\add_35/carry[1] ), 
        .CO(\add_35/carry[2] ), .S(q_res[1]) );
  FA_X1 \add_35/U1_2  ( .A(N2), .B(warp_num_in[2]), .CI(\add_35/carry[2] ), 
        .CO(\add_35/carry[3] ), .S(q_res[2]) );
  FA_X1 \add_35/U1_3  ( .A(N3), .B(warp_num_in[3]), .CI(\add_35/carry[3] ), 
        .CO(\add_35/carry[4] ), .S(q_res[3]) );
  FA_X1 \add_35/U1_4  ( .A(N4), .B(warp_num_in[4]), .CI(\add_35/carry[4] ), 
        .CO(\add_35/carry[5] ), .S(q_res[4]) );
  XOR2_X1 U3 ( .A(N9), .B(\add_35/carry[9] ), .Z(q_res[9]) );
  AND2_X1 U4 ( .A1(N8), .A2(\add_35/carry[8] ), .ZN(\add_35/carry[9] ) );
  XOR2_X1 U5 ( .A(N8), .B(\add_35/carry[8] ), .Z(q_res[8]) );
  AND2_X1 U6 ( .A1(N7), .A2(\add_35/carry[7] ), .ZN(\add_35/carry[8] ) );
  XOR2_X1 U7 ( .A(N7), .B(\add_35/carry[7] ), .Z(q_res[7]) );
  AND2_X1 U8 ( .A1(N6), .A2(\add_35/carry[6] ), .ZN(\add_35/carry[7] ) );
  XOR2_X1 U9 ( .A(N6), .B(\add_35/carry[6] ), .Z(q_res[6]) );
  AND2_X1 U10 ( .A1(N5), .A2(\add_35/carry[5] ), .ZN(\add_35/carry[6] ) );
  XOR2_X1 U11 ( .A(N5), .B(\add_35/carry[5] ), .Z(q_res[5]) );
  AND2_X1 U12 ( .A1(warp_num_in[0]), .A2(N0), .ZN(\add_35/carry[1] ) );
  XOR2_X1 U13 ( .A(warp_num_in[0]), .B(N0), .Z(warp_id_out[0]) );
  MUX2_X1 U14 ( .A(q_res[1]), .B(q_res[1]), .S(\rem_36/u_div/PartRem[1><5] ), 
        .Z(warp_id_out[1]) );
  MUX2_X1 U15 ( .A(q_res[2]), .B(q_res[2]), .S(\rem_36/u_div/PartRem[2><5] ), 
        .Z(\rem_36/u_div/PartRem[1><2] ) );
  MUX2_X1 U16 ( .A(\rem_36/u_div/PartRem[1><2] ), .B(
        \rem_36/u_div/PartRem[1><2] ), .S(\rem_36/u_div/PartRem[1><5] ), .Z(
        warp_id_out[2]) );
  MUX2_X1 U17 ( .A(q_res[3]), .B(q_res[3]), .S(\rem_36/u_div/PartRem[3><5] ), 
        .Z(\rem_36/u_div/PartRem[2><2] ) );
  MUX2_X1 U18 ( .A(\rem_36/u_div/PartRem[2><2] ), .B(
        \rem_36/u_div/PartRem[2><2] ), .S(\rem_36/u_div/PartRem[2><5] ), .Z(
        \rem_36/u_div/PartRem[1><3] ) );
  MUX2_X1 U19 ( .A(\rem_36/u_div/PartRem[1><3] ), .B(
        \rem_36/u_div/PartRem[1><3] ), .S(\rem_36/u_div/PartRem[1><5] ), .Z(
        warp_id_out[3]) );
  MUX2_X1 U20 ( .A(q_res[4]), .B(q_res[4]), .S(\rem_36/u_div/PartRem[4><5] ), 
        .Z(\rem_36/u_div/PartRem[3><2] ) );
  MUX2_X1 U21 ( .A(\rem_36/u_div/PartRem[3><2] ), .B(
        \rem_36/u_div/PartRem[3><2] ), .S(\rem_36/u_div/PartRem[3><5] ), .Z(
        \rem_36/u_div/PartRem[2><3] ) );
  MUX2_X1 U22 ( .A(\rem_36/u_div/PartRem[2><3] ), .B(
        \rem_36/u_div/PartRem[2><3] ), .S(\rem_36/u_div/PartRem[2><5] ), .Z(
        \rem_36/u_div/PartRem[1><4] ) );
  MUX2_X1 U23 ( .A(\rem_36/u_div/PartRem[1><4] ), .B(
        \rem_36/u_div/PartRem[1><4] ), .S(\rem_36/u_div/PartRem[1><5] ), .Z(
        warp_id_out[4]) );
  MUX2_X1 U24 ( .A(q_res[5]), .B(q_res[5]), .S(q_res[9]), .Z(
        \rem_36/u_div/PartRem[4><2] ) );
  MUX2_X1 U25 ( .A(\rem_36/u_div/PartRem[4><2] ), .B(
        \rem_36/u_div/PartRem[4><2] ), .S(\rem_36/u_div/PartRem[4><5] ), .Z(
        \rem_36/u_div/PartRem[3><3] ) );
  MUX2_X1 U26 ( .A(\rem_36/u_div/PartRem[3><3] ), .B(
        \rem_36/u_div/PartRem[3><3] ), .S(\rem_36/u_div/PartRem[3><5] ), .Z(
        \rem_36/u_div/PartRem[2><4] ) );
  MUX2_X1 U27 ( .A(\rem_36/u_div/PartRem[2><4] ), .B(
        \rem_36/u_div/PartRem[2><4] ), .S(\rem_36/u_div/PartRem[2><5] ), .Z(
        \rem_36/u_div/PartRem[1><5] ) );
  MUX2_X1 U28 ( .A(q_res[6]), .B(q_res[6]), .S(q_res[9]), .Z(
        \rem_36/u_div/PartRem[4><3] ) );
  MUX2_X1 U29 ( .A(\rem_36/u_div/PartRem[4><3] ), .B(
        \rem_36/u_div/PartRem[4><3] ), .S(\rem_36/u_div/PartRem[4><5] ), .Z(
        \rem_36/u_div/PartRem[3><4] ) );
  MUX2_X1 U30 ( .A(\rem_36/u_div/PartRem[3><4] ), .B(
        \rem_36/u_div/PartRem[3><4] ), .S(\rem_36/u_div/PartRem[3><5] ), .Z(
        \rem_36/u_div/PartRem[2><5] ) );
  MUX2_X1 U31 ( .A(q_res[7]), .B(q_res[7]), .S(q_res[9]), .Z(
        \rem_36/u_div/PartRem[4><4] ) );
  MUX2_X1 U32 ( .A(\rem_36/u_div/PartRem[4><4] ), .B(
        \rem_36/u_div/PartRem[4><4] ), .S(\rem_36/u_div/PartRem[4><5] ), .Z(
        \rem_36/u_div/PartRem[3><5] ) );
  MUX2_X1 U33 ( .A(q_res[8]), .B(q_res[8]), .S(q_res[9]), .Z(
        \rem_36/u_div/PartRem[4><5] ) );
endmodule

/* -------------------------------------------------------------------------
-- Company:          
-- Engineer:         
-- 
-- Create Date:      
-- Module Name:      warp_scheduler - post_syn. 
-- Project Name:     GPGPU
-- Target Devices: 
-- Tool versions:    
-- Description: 
--
----------------------------------------------------------------------------
---------------------------------------------------------------------------- */

module warp_scheduler_SHMEM_ADDR_SIZE14_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, 
        GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  INV_X1 U1 ( .A(A[1]), .ZN(n2) );
  INV_X1 U2 ( .A(A[0]), .ZN(n3) );
  INV_X1 U3 ( .A(B[1]), .ZN(n1) );
  NOR4_X1 U4 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(EQ) );
  NAND4_X1 U5 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .ZN(n7) );
  XNOR2_X1 U6 ( .A(B[3]), .B(A[3]), .ZN(n11) );
  XNOR2_X1 U7 ( .A(B[4]), .B(A[4]), .ZN(n10) );
  XNOR2_X1 U8 ( .A(B[5]), .B(A[5]), .ZN(n9) );
  XNOR2_X1 U9 ( .A(B[6]), .B(A[6]), .ZN(n8) );
  NAND4_X1 U10 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .ZN(n6) );
  OAI22_X1 U11 ( .A1(n16), .A2(n2), .B1(B[1]), .B2(n16), .ZN(n15) );
  AND2_X1 U12 ( .A1(B[0]), .A2(n3), .ZN(n16) );
  OAI22_X1 U13 ( .A1(A[1]), .A2(n17), .B1(n17), .B2(n1), .ZN(n14) );
  NOR2_X1 U14 ( .A1(n3), .A2(B[0]), .ZN(n17) );
  XNOR2_X1 U15 ( .A(B[31]), .B(A[31]), .ZN(n13) );
  XNOR2_X1 U16 ( .A(B[2]), .B(A[2]), .ZN(n12) );
  NAND2_X1 U17 ( .A1(n18), .A2(n19), .ZN(n5) );
  NOR4_X1 U18 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n19) );
  XOR2_X1 U19 ( .A(B[10]), .B(A[10]), .Z(n23) );
  XOR2_X1 U20 ( .A(B[9]), .B(A[9]), .Z(n22) );
  XOR2_X1 U21 ( .A(B[8]), .B(A[8]), .Z(n21) );
  XOR2_X1 U22 ( .A(B[7]), .B(A[7]), .Z(n20) );
  NOR4_X1 U23 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n18) );
  XOR2_X1 U24 ( .A(B[14]), .B(A[14]), .Z(n27) );
  XOR2_X1 U25 ( .A(B[13]), .B(A[13]), .Z(n26) );
  XOR2_X1 U26 ( .A(B[12]), .B(A[12]), .Z(n25) );
  XOR2_X1 U27 ( .A(B[11]), .B(A[11]), .Z(n24) );
  NAND4_X1 U28 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n4) );
  NOR4_X1 U29 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(n31) );
  XOR2_X1 U30 ( .A(B[18]), .B(A[18]), .Z(n35) );
  XOR2_X1 U31 ( .A(B[17]), .B(A[17]), .Z(n34) );
  XOR2_X1 U32 ( .A(B[16]), .B(A[16]), .Z(n33) );
  XOR2_X1 U33 ( .A(B[15]), .B(A[15]), .Z(n32) );
  NOR4_X1 U34 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n30) );
  XOR2_X1 U35 ( .A(B[22]), .B(A[22]), .Z(n39) );
  XOR2_X1 U36 ( .A(B[21]), .B(A[21]), .Z(n38) );
  XOR2_X1 U37 ( .A(B[20]), .B(A[20]), .Z(n37) );
  XOR2_X1 U38 ( .A(B[19]), .B(A[19]), .Z(n36) );
  NOR4_X1 U39 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n29) );
  XOR2_X1 U40 ( .A(B[26]), .B(A[26]), .Z(n43) );
  XOR2_X1 U41 ( .A(B[25]), .B(A[25]), .Z(n42) );
  XOR2_X1 U42 ( .A(B[24]), .B(A[24]), .Z(n41) );
  XOR2_X1 U43 ( .A(B[23]), .B(A[23]), .Z(n40) );
  NOR4_X1 U44 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n28) );
  XOR2_X1 U45 ( .A(B[30]), .B(A[30]), .Z(n47) );
  XOR2_X1 U46 ( .A(B[29]), .B(A[29]), .Z(n46) );
  XOR2_X1 U47 ( .A(B[28]), .B(A[28]), .Z(n45) );
  XOR2_X1 U48 ( .A(B[27]), .B(A[27]), .Z(n44) );
endmodule



module warp_scheduler ( clk_in, host_reset, reset, 
        pipeline_stall_in, num_blocks_in, num_warps_in, gprs_size_in, 
        warps_done_mask_in, warp_pool_addr_out, warp_pool_wr_en_out, 
        warp_pool_wr_data_out, warp_pool_rd_data_in, warp_state_addr_out, 
        warp_state_wr_en_out, warp_state_wr_data_out, warp_state_rd_data_in, 
        program_cntr_out, warp_id_out, warp_lane_id_out, cta_id_out, 
        initial_mask_out, current_mask_out, shmem_base_addr_out, gprs_size_out, 
        gprs_base_addr_out, done, pipeline_warpunit_done, fetch_en );
  input [3:0] num_blocks_in;
  input [4:0] num_warps_in;
  input [8:0] gprs_size_in;
  input [31:0] warps_done_mask_in;
  output [4:0] warp_pool_addr_out;
  output [127:0] warp_pool_wr_data_out;
  input [127:0] warp_pool_rd_data_in;
  output [4:0] warp_state_addr_out;
  output [1:0] warp_state_wr_data_out;
  input [1:0] warp_state_rd_data_in;
  output [31:0] program_cntr_out;
  output [4:0] warp_id_out;
  output [1:0] warp_lane_id_out;
  output [3:0] cta_id_out;
  output [31:0] initial_mask_out;
  output [31:0] current_mask_out;
  output [13:0] shmem_base_addr_out;
  output [8:0] gprs_size_out;
  output [8:0] gprs_base_addr_out;
  input clk_in, host_reset, reset, pipeline_stall_in;
  output warp_pool_wr_en_out, warp_state_wr_en_out, done,
         pipeline_warpunit_done, fetch_en;
  wire   N52, N63, N64, N66, N67, N70, N71, N72, N73, N94, N321, N322, N323,
         N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334,
         N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345,
         N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356,
         N357, N358, N359, N360, N362, N364, N365, N366, N367, N368, N369,
         N370, N371, N372, N373, N375, N376, N377, N378, N379, N380, N381,
         N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392,
         N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403,
         N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414,
         N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425,
         N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436,
         N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447,
         N448, N449, N450, N451, N452, N453, N454, N455, n161, n166, n167,
         n168, n169, n170, n177, n178, n179, n180, n181, n182, n183, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         \r149/carry[4] , \r149/carry[3] , \r149/carry[2] , n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n162, n163, n164, n165, n171,
         n172, n173, n174, n175, n176, n184, n185, n186, n187, n212, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649;
  wire   [1:0] warp_lane_cnt;
  wire   [4:0] warp_id_cnt;
  wire   [2:0] warp_scheduler_next_state;
  wire   [2:0] warp_scheduler_state_machine;
  wire   [31:0] warps_done_mask;
  assign warp_pool_wr_en_out = 1'b0;
  assign warp_state_wr_data_out[1] = 1'b0;
  assign N321 = warp_pool_rd_data_in[110];
  assign N322 = warp_pool_rd_data_in[111];
  assign N323 = warp_pool_rd_data_in[112];
  assign N324 = warp_pool_rd_data_in[113];
  assign N325 = warp_pool_rd_data_in[114];
  assign N326 = warp_pool_rd_data_in[115];
  assign N327 = warp_pool_rd_data_in[116];
  assign N328 = warp_pool_rd_data_in[117];
  assign N329 = warp_pool_rd_data_in[118];
  assign N330 = warp_pool_rd_data_in[119];
  assign N331 = warp_pool_rd_data_in[120];
  assign N332 = warp_pool_rd_data_in[121];
  assign N333 = warp_pool_rd_data_in[122];
  assign N334 = warp_pool_rd_data_in[123];
  assign N335 = warp_pool_rd_data_in[106];
  assign N336 = warp_pool_rd_data_in[107];
  assign N337 = warp_pool_rd_data_in[108];
  assign N338 = warp_pool_rd_data_in[109];
  assign N339 = warp_pool_rd_data_in[97];
  assign N340 = warp_pool_rd_data_in[98];
  assign N341 = warp_pool_rd_data_in[99];
  assign N342 = warp_pool_rd_data_in[100];
  assign N343 = warp_pool_rd_data_in[101];
  assign N344 = warp_pool_rd_data_in[102];
  assign N345 = warp_pool_rd_data_in[103];
  assign N346 = warp_pool_rd_data_in[104];
  assign N347 = warp_pool_rd_data_in[105];
  assign N348 = warp_pool_rd_data_in[32];
  assign N349 = warp_pool_rd_data_in[33];
  assign N350 = warp_pool_rd_data_in[34];
  assign N351 = warp_pool_rd_data_in[35];
  assign N352 = warp_pool_rd_data_in[36];
  assign N353 = warp_pool_rd_data_in[37];
  assign N354 = warp_pool_rd_data_in[38];
  assign N355 = warp_pool_rd_data_in[39];
  assign N356 = warp_pool_rd_data_in[40];
  assign N357 = warp_pool_rd_data_in[41];
  assign N358 = warp_pool_rd_data_in[42];
  assign N359 = warp_pool_rd_data_in[43];
  assign N360 = warp_pool_rd_data_in[44];
  assign N362 = warp_pool_rd_data_in[45];
  assign N364 = warp_pool_rd_data_in[46];
  assign N365 = warp_pool_rd_data_in[47];
  assign N366 = warp_pool_rd_data_in[48];
  assign N367 = warp_pool_rd_data_in[49];
  assign N368 = warp_pool_rd_data_in[50];
  assign N369 = warp_pool_rd_data_in[51];
  assign N370 = warp_pool_rd_data_in[52];
  assign N371 = warp_pool_rd_data_in[53];
  assign N372 = warp_pool_rd_data_in[54];
  assign N373 = warp_pool_rd_data_in[55];
  assign N375 = warp_pool_rd_data_in[56];
  assign N376 = warp_pool_rd_data_in[57];
  assign N377 = warp_pool_rd_data_in[58];
  assign N378 = warp_pool_rd_data_in[59];
  assign N379 = warp_pool_rd_data_in[60];
  assign N380 = warp_pool_rd_data_in[61];
  assign N381 = warp_pool_rd_data_in[62];
  assign N382 = warp_pool_rd_data_in[63];
  assign N383 = warp_pool_rd_data_in[0];
  assign N384 = warp_pool_rd_data_in[1];
  assign N385 = warp_pool_rd_data_in[2];
  assign N386 = warp_pool_rd_data_in[3];
  assign N387 = warp_pool_rd_data_in[4];
  assign N388 = warp_pool_rd_data_in[5];
  assign N389 = warp_pool_rd_data_in[6];
  assign N390 = warp_pool_rd_data_in[7];
  assign N391 = warp_pool_rd_data_in[8];
  assign N392 = warp_pool_rd_data_in[9];
  assign N393 = warp_pool_rd_data_in[10];
  assign N394 = warp_pool_rd_data_in[11];
  assign N395 = warp_pool_rd_data_in[12];
  assign N396 = warp_pool_rd_data_in[13];
  assign N397 = warp_pool_rd_data_in[14];
  assign N398 = warp_pool_rd_data_in[15];
  assign N399 = warp_pool_rd_data_in[16];
  assign N400 = warp_pool_rd_data_in[17];
  assign N401 = warp_pool_rd_data_in[18];
  assign N402 = warp_pool_rd_data_in[19];
  assign N403 = warp_pool_rd_data_in[20];
  assign N404 = warp_pool_rd_data_in[21];
  assign N405 = warp_pool_rd_data_in[22];
  assign N406 = warp_pool_rd_data_in[23];
  assign N407 = warp_pool_rd_data_in[24];
  assign N408 = warp_pool_rd_data_in[25];
  assign N409 = warp_pool_rd_data_in[26];
  assign N410 = warp_pool_rd_data_in[27];
  assign N411 = warp_pool_rd_data_in[28];
  assign N412 = warp_pool_rd_data_in[29];
  assign N413 = warp_pool_rd_data_in[30];
  assign N414 = warp_pool_rd_data_in[31];
  assign N415 = warp_pool_rd_data_in[64];
  assign N416 = warp_pool_rd_data_in[65];
  assign N417 = warp_pool_rd_data_in[66];
  assign N418 = warp_pool_rd_data_in[67];
  assign N419 = warp_pool_rd_data_in[68];
  assign N420 = warp_pool_rd_data_in[69];
  assign N421 = warp_pool_rd_data_in[70];
  assign N422 = warp_pool_rd_data_in[71];
  assign N423 = warp_pool_rd_data_in[72];
  assign N424 = warp_pool_rd_data_in[73];
  assign N425 = warp_pool_rd_data_in[74];
  assign N426 = warp_pool_rd_data_in[75];
  assign N427 = warp_pool_rd_data_in[76];
  assign N428 = warp_pool_rd_data_in[77];
  assign N429 = warp_pool_rd_data_in[78];
  assign N430 = warp_pool_rd_data_in[79];
  assign N431 = warp_pool_rd_data_in[80];
  assign N432 = warp_pool_rd_data_in[81];
  assign N433 = warp_pool_rd_data_in[82];
  assign N434 = warp_pool_rd_data_in[83];
  assign N435 = warp_pool_rd_data_in[84];
  assign N436 = warp_pool_rd_data_in[85];
  assign N437 = warp_pool_rd_data_in[86];
  assign N438 = warp_pool_rd_data_in[87];
  assign N439 = warp_pool_rd_data_in[88];
  assign N440 = warp_pool_rd_data_in[89];
  assign N441 = warp_pool_rd_data_in[90];
  assign N442 = warp_pool_rd_data_in[91];
  assign N443 = warp_pool_rd_data_in[92];
  assign N444 = warp_pool_rd_data_in[93];
  assign N445 = warp_pool_rd_data_in[94];
  assign N446 = warp_pool_rd_data_in[95];
  assign N447 = gprs_size_in[0];
  assign N448 = gprs_size_in[1];
  assign N449 = gprs_size_in[2];
  assign N450 = gprs_size_in[3];
  assign N451 = gprs_size_in[4];
  assign N452 = gprs_size_in[5];
  assign N453 = gprs_size_in[6];
  assign N454 = gprs_size_in[7];
  assign N455 = gprs_size_in[8];
  assign warp_pool_wr_data_out[127] = 1'b0;
  assign warp_pool_wr_data_out[126] = 1'b0;
  assign warp_pool_wr_data_out[125] = 1'b0;
  assign warp_pool_wr_data_out[124] = 1'b0;
  assign warp_pool_wr_data_out[123] = 1'b0;
  assign warp_pool_wr_data_out[122] = 1'b0;
  assign warp_pool_wr_data_out[121] = 1'b0;
  assign warp_pool_wr_data_out[120] = 1'b0;
  assign warp_pool_wr_data_out[119] = 1'b0;
  assign warp_pool_wr_data_out[118] = 1'b0;
  assign warp_pool_wr_data_out[117] = 1'b0;
  assign warp_pool_wr_data_out[116] = 1'b0;
  assign warp_pool_wr_data_out[115] = 1'b0;
  assign warp_pool_wr_data_out[114] = 1'b0;
  assign warp_pool_wr_data_out[113] = 1'b0;
  assign warp_pool_wr_data_out[112] = 1'b0;
  assign warp_pool_wr_data_out[111] = 1'b0;
  assign warp_pool_wr_data_out[110] = 1'b0;
  assign warp_pool_wr_data_out[109] = 1'b0;
  assign warp_pool_wr_data_out[108] = 1'b0;
  assign warp_pool_wr_data_out[107] = 1'b0;
  assign warp_pool_wr_data_out[106] = 1'b0;
  assign warp_pool_wr_data_out[105] = 1'b0;
  assign warp_pool_wr_data_out[104] = 1'b0;
  assign warp_pool_wr_data_out[103] = 1'b0;
  assign warp_pool_wr_data_out[102] = 1'b0;
  assign warp_pool_wr_data_out[101] = 1'b0;
  assign warp_pool_wr_data_out[100] = 1'b0;
  assign warp_pool_wr_data_out[99] = 1'b0;
  assign warp_pool_wr_data_out[98] = 1'b0;
  assign warp_pool_wr_data_out[97] = 1'b0;
  assign warp_pool_wr_data_out[96] = 1'b0;
  assign warp_pool_wr_data_out[95] = 1'b0;
  assign warp_pool_wr_data_out[94] = 1'b0;
  assign warp_pool_wr_data_out[93] = 1'b0;
  assign warp_pool_wr_data_out[92] = 1'b0;
  assign warp_pool_wr_data_out[91] = 1'b0;
  assign warp_pool_wr_data_out[90] = 1'b0;
  assign warp_pool_wr_data_out[89] = 1'b0;
  assign warp_pool_wr_data_out[88] = 1'b0;
  assign warp_pool_wr_data_out[87] = 1'b0;
  assign warp_pool_wr_data_out[86] = 1'b0;
  assign warp_pool_wr_data_out[85] = 1'b0;
  assign warp_pool_wr_data_out[84] = 1'b0;
  assign warp_pool_wr_data_out[83] = 1'b0;
  assign warp_pool_wr_data_out[82] = 1'b0;
  assign warp_pool_wr_data_out[81] = 1'b0;
  assign warp_pool_wr_data_out[80] = 1'b0;
  assign warp_pool_wr_data_out[79] = 1'b0;
  assign warp_pool_wr_data_out[78] = 1'b0;
  assign warp_pool_wr_data_out[77] = 1'b0;
  assign warp_pool_wr_data_out[76] = 1'b0;
  assign warp_pool_wr_data_out[75] = 1'b0;
  assign warp_pool_wr_data_out[74] = 1'b0;
  assign warp_pool_wr_data_out[73] = 1'b0;
  assign warp_pool_wr_data_out[72] = 1'b0;
  assign warp_pool_wr_data_out[71] = 1'b0;
  assign warp_pool_wr_data_out[70] = 1'b0;
  assign warp_pool_wr_data_out[69] = 1'b0;
  assign warp_pool_wr_data_out[68] = 1'b0;
  assign warp_pool_wr_data_out[67] = 1'b0;
  assign warp_pool_wr_data_out[66] = 1'b0;
  assign warp_pool_wr_data_out[65] = 1'b0;
  assign warp_pool_wr_data_out[64] = 1'b0;
  assign warp_pool_wr_data_out[63] = 1'b0;
  assign warp_pool_wr_data_out[62] = 1'b0;
  assign warp_pool_wr_data_out[61] = 1'b0;
  assign warp_pool_wr_data_out[60] = 1'b0;
  assign warp_pool_wr_data_out[59] = 1'b0;
  assign warp_pool_wr_data_out[58] = 1'b0;
  assign warp_pool_wr_data_out[57] = 1'b0;
  assign warp_pool_wr_data_out[56] = 1'b0;
  assign warp_pool_wr_data_out[55] = 1'b0;
  assign warp_pool_wr_data_out[54] = 1'b0;
  assign warp_pool_wr_data_out[53] = 1'b0;
  assign warp_pool_wr_data_out[52] = 1'b0;
  assign warp_pool_wr_data_out[51] = 1'b0;
  assign warp_pool_wr_data_out[50] = 1'b0;
  assign warp_pool_wr_data_out[49] = 1'b0;
  assign warp_pool_wr_data_out[48] = 1'b0;
  assign warp_pool_wr_data_out[47] = 1'b0;
  assign warp_pool_wr_data_out[46] = 1'b0;
  assign warp_pool_wr_data_out[45] = 1'b0;
  assign warp_pool_wr_data_out[44] = 1'b0;
  assign warp_pool_wr_data_out[43] = 1'b0;
  assign warp_pool_wr_data_out[42] = 1'b0;
  assign warp_pool_wr_data_out[41] = 1'b0;
  assign warp_pool_wr_data_out[40] = 1'b0;
  assign warp_pool_wr_data_out[39] = 1'b0;
  assign warp_pool_wr_data_out[38] = 1'b0;
  assign warp_pool_wr_data_out[37] = 1'b0;
  assign warp_pool_wr_data_out[36] = 1'b0;
  assign warp_pool_wr_data_out[35] = 1'b0;
  assign warp_pool_wr_data_out[34] = 1'b0;
  assign warp_pool_wr_data_out[33] = 1'b0;
  assign warp_pool_wr_data_out[32] = 1'b0;
  assign warp_pool_wr_data_out[31] = 1'b0;
  assign warp_pool_wr_data_out[30] = 1'b0;
  assign warp_pool_wr_data_out[29] = 1'b0;
  assign warp_pool_wr_data_out[28] = 1'b0;
  assign warp_pool_wr_data_out[27] = 1'b0;
  assign warp_pool_wr_data_out[26] = 1'b0;
  assign warp_pool_wr_data_out[25] = 1'b0;
  assign warp_pool_wr_data_out[24] = 1'b0;
  assign warp_pool_wr_data_out[23] = 1'b0;
  assign warp_pool_wr_data_out[22] = 1'b0;
  assign warp_pool_wr_data_out[21] = 1'b0;
  assign warp_pool_wr_data_out[20] = 1'b0;
  assign warp_pool_wr_data_out[19] = 1'b0;
  assign warp_pool_wr_data_out[18] = 1'b0;
  assign warp_pool_wr_data_out[17] = 1'b0;
  assign warp_pool_wr_data_out[16] = 1'b0;
  assign warp_pool_wr_data_out[15] = 1'b0;
  assign warp_pool_wr_data_out[14] = 1'b0;
  assign warp_pool_wr_data_out[13] = 1'b0;
  assign warp_pool_wr_data_out[12] = 1'b0;
  assign warp_pool_wr_data_out[11] = 1'b0;
  assign warp_pool_wr_data_out[10] = 1'b0;
  assign warp_pool_wr_data_out[9] = 1'b0;
  assign warp_pool_wr_data_out[8] = 1'b0;
  assign warp_pool_wr_data_out[7] = 1'b0;
  assign warp_pool_wr_data_out[6] = 1'b0;
  assign warp_pool_wr_data_out[5] = 1'b0;
  assign warp_pool_wr_data_out[4] = 1'b0;
  assign warp_pool_wr_data_out[3] = 1'b0;
  assign warp_pool_wr_data_out[2] = 1'b0;
  assign warp_pool_wr_data_out[1] = 1'b0;
  assign warp_pool_wr_data_out[0] = 1'b0;

  DFFR_X1 \warp_scheduler_next_state_reg[0]  ( .D(n430), .CK(clk_in), .RN(n150), .Q(warp_scheduler_next_state[0]), .QN(n183) );
  DFFR_X1 \warp_scheduler_state_machine_reg[0]  ( .D(n428), .CK(clk_in), .RN(
        n150), .Q(warp_scheduler_state_machine[0]), .QN(n167) );
  DFFR_X1 \warp_lane_cnt_reg[1]  ( .D(n425), .CK(clk_in), .RN(n150), .Q(
        warp_lane_cnt[1]), .QN(n168) );
  DFFR_X1 \warp_scheduler_next_state_reg[2]  ( .D(n421), .CK(clk_in), .RN(n150), .Q(warp_scheduler_next_state[2]), .QN(n181) );
  DFFR_X1 \warp_scheduler_state_machine_reg[2]  ( .D(n429), .CK(clk_in), .RN(
        n150), .Q(warp_scheduler_state_machine[2]), .QN(n161) );
  DFFR_X1 \initial_mask_out_reg[12]  ( .D(n500), .CK(clk_in), .RN(n150), .Q(
        initial_mask_out[12]) );
  DFFR_X1 \initial_mask_out_reg[11]  ( .D(n501), .CK(clk_in), .RN(n150), .Q(
        initial_mask_out[11]) );
  DFFR_X1 \initial_mask_out_reg[10]  ( .D(n502), .CK(clk_in), .RN(n150), .Q(
        initial_mask_out[10]) );
  DFFR_X1 \initial_mask_out_reg[9]  ( .D(n503), .CK(clk_in), .RN(n150), .Q(
        initial_mask_out[9]) );
  DFFR_X1 \initial_mask_out_reg[8]  ( .D(n504), .CK(clk_in), .RN(n150), .Q(
        initial_mask_out[8]) );
  DFFR_X1 \initial_mask_out_reg[7]  ( .D(n505), .CK(clk_in), .RN(n150), .Q(
        initial_mask_out[7]) );
  DFFR_X1 \initial_mask_out_reg[6]  ( .D(n506), .CK(clk_in), .RN(n149), .Q(
        initial_mask_out[6]) );
  DFFR_X1 \initial_mask_out_reg[5]  ( .D(n507), .CK(clk_in), .RN(n149), .Q(
        initial_mask_out[5]) );
  DFFR_X1 \initial_mask_out_reg[4]  ( .D(n508), .CK(clk_in), .RN(n149), .Q(
        initial_mask_out[4]) );
  DFFR_X1 \initial_mask_out_reg[3]  ( .D(n509), .CK(clk_in), .RN(n149), .Q(
        initial_mask_out[3]) );
  DFFR_X1 \initial_mask_out_reg[2]  ( .D(n510), .CK(clk_in), .RN(n149), .Q(
        initial_mask_out[2]) );
  DFFR_X1 \initial_mask_out_reg[1]  ( .D(n511), .CK(clk_in), .RN(n149), .Q(
        initial_mask_out[1]) );
  DFFR_X1 \initial_mask_out_reg[0]  ( .D(n512), .CK(clk_in), .RN(n149), .Q(
        initial_mask_out[0]) );
  DFFR_X1 \gprs_base_addr_out_reg[8]  ( .D(n513), .CK(clk_in), .RN(n149), .Q(
        gprs_base_addr_out[8]) );
  DFFR_X1 \gprs_base_addr_out_reg[7]  ( .D(n514), .CK(clk_in), .RN(n149), .Q(
        gprs_base_addr_out[7]) );
  DFFR_X1 \gprs_base_addr_out_reg[6]  ( .D(n515), .CK(clk_in), .RN(n149), .Q(
        gprs_base_addr_out[6]) );
  DFFR_X1 \gprs_base_addr_out_reg[5]  ( .D(n516), .CK(clk_in), .RN(n149), .Q(
        gprs_base_addr_out[5]) );
  DFFR_X1 \gprs_base_addr_out_reg[4]  ( .D(n517), .CK(clk_in), .RN(n149), .Q(
        gprs_base_addr_out[4]) );
  DFFR_X1 \gprs_base_addr_out_reg[3]  ( .D(n518), .CK(clk_in), .RN(n148), .Q(
        gprs_base_addr_out[3]) );
  DFFR_X1 \gprs_base_addr_out_reg[2]  ( .D(n519), .CK(clk_in), .RN(n148), .Q(
        gprs_base_addr_out[2]) );
  DFFR_X1 \gprs_base_addr_out_reg[1]  ( .D(n520), .CK(clk_in), .RN(n148), .Q(
        gprs_base_addr_out[1]) );
  DFFR_X1 \gprs_base_addr_out_reg[0]  ( .D(n521), .CK(clk_in), .RN(n148), .Q(
        gprs_base_addr_out[0]) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n522), .CK(clk_in), .RN(n148), .Q(
        cta_id_out[3]) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n523), .CK(clk_in), .RN(n148), .Q(
        cta_id_out[2]) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n524), .CK(clk_in), .RN(n148), .Q(
        cta_id_out[1]) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n525), .CK(clk_in), .RN(n148), .Q(
        cta_id_out[0]) );
  DFFR_X1 \shmem_base_addr_out_reg[13]  ( .D(n526), .CK(clk_in), .RN(n148), 
        .Q(shmem_base_addr_out[13]) );
  DFFR_X1 \shmem_base_addr_out_reg[12]  ( .D(n527), .CK(clk_in), .RN(n148), 
        .Q(shmem_base_addr_out[12]) );
  DFFR_X1 \shmem_base_addr_out_reg[11]  ( .D(n528), .CK(clk_in), .RN(n148), 
        .Q(shmem_base_addr_out[11]) );
  DFFR_X1 \shmem_base_addr_out_reg[10]  ( .D(n529), .CK(clk_in), .RN(n148), 
        .Q(shmem_base_addr_out[10]) );
  DFFR_X1 \shmem_base_addr_out_reg[9]  ( .D(n530), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[9]) );
  DFFR_X1 \shmem_base_addr_out_reg[8]  ( .D(n531), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[8]) );
  DFFR_X1 \shmem_base_addr_out_reg[7]  ( .D(n532), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[7]) );
  DFFR_X1 \shmem_base_addr_out_reg[6]  ( .D(n533), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[6]) );
  DFFR_X1 \shmem_base_addr_out_reg[5]  ( .D(n534), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[5]) );
  DFFR_X1 \shmem_base_addr_out_reg[4]  ( .D(n535), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[4]) );
  DFFR_X1 \shmem_base_addr_out_reg[3]  ( .D(n536), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[3]) );
  DFFR_X1 \shmem_base_addr_out_reg[2]  ( .D(n537), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[2]) );
  DFFR_X1 \shmem_base_addr_out_reg[1]  ( .D(n538), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[1]) );
  DFFR_X1 \shmem_base_addr_out_reg[0]  ( .D(n539), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[0]) );
  DFFR_X1 \gprs_size_out_reg[8]  ( .D(n540), .CK(clk_in), .RN(n147), .Q(
        gprs_size_out[8]) );
  DFFR_X1 \gprs_size_out_reg[7]  ( .D(n541), .CK(clk_in), .RN(n147), .Q(
        gprs_size_out[7]) );
  DFFR_X1 \gprs_size_out_reg[6]  ( .D(n542), .CK(clk_in), .RN(n146), .Q(
        gprs_size_out[6]) );
  DFFR_X1 \gprs_size_out_reg[5]  ( .D(n543), .CK(clk_in), .RN(n146), .Q(
        gprs_size_out[5]) );
  DFFR_X1 \gprs_size_out_reg[4]  ( .D(n544), .CK(clk_in), .RN(n146), .Q(
        gprs_size_out[4]) );
  DFFR_X1 \gprs_size_out_reg[3]  ( .D(n545), .CK(clk_in), .RN(n146), .Q(
        gprs_size_out[3]) );
  DFFR_X1 \gprs_size_out_reg[2]  ( .D(n546), .CK(clk_in), .RN(n146), .Q(
        gprs_size_out[2]) );
  DFFR_X1 \gprs_size_out_reg[1]  ( .D(n547), .CK(clk_in), .RN(n146), .Q(
        gprs_size_out[1]) );
  DFFR_X1 \gprs_size_out_reg[0]  ( .D(n548), .CK(clk_in), .RN(n146), .Q(
        gprs_size_out[0]) );
  DFFR_X1 \program_cntr_out_reg[31]  ( .D(n549), .CK(clk_in), .RN(n146), .Q(
        program_cntr_out[31]) );
  DFFR_X1 \program_cntr_out_reg[30]  ( .D(n550), .CK(clk_in), .RN(n146), .Q(
        program_cntr_out[30]) );
  DFFR_X1 \program_cntr_out_reg[29]  ( .D(n551), .CK(clk_in), .RN(n146), .Q(
        program_cntr_out[29]) );
  DFFR_X1 \program_cntr_out_reg[28]  ( .D(n552), .CK(clk_in), .RN(n146), .Q(
        program_cntr_out[28]) );
  DFFR_X1 \program_cntr_out_reg[27]  ( .D(n553), .CK(clk_in), .RN(n146), .Q(
        program_cntr_out[27]) );
  DFFR_X1 \program_cntr_out_reg[26]  ( .D(n554), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[26]) );
  DFFR_X1 \program_cntr_out_reg[25]  ( .D(n555), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[25]) );
  DFFR_X1 \program_cntr_out_reg[24]  ( .D(n556), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[24]) );
  DFFR_X1 \program_cntr_out_reg[23]  ( .D(n557), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[23]) );
  DFFR_X1 \program_cntr_out_reg[22]  ( .D(n558), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[22]) );
  DFFR_X1 \program_cntr_out_reg[21]  ( .D(n559), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[21]) );
  DFFR_X1 \program_cntr_out_reg[20]  ( .D(n560), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[20]) );
  DFFR_X1 \program_cntr_out_reg[19]  ( .D(n561), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[19]) );
  DFFR_X1 \program_cntr_out_reg[18]  ( .D(n562), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[18]) );
  DFFR_X1 \program_cntr_out_reg[17]  ( .D(n563), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[17]) );
  DFFR_X1 \program_cntr_out_reg[16]  ( .D(n564), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[16]) );
  DFFR_X1 \program_cntr_out_reg[15]  ( .D(n565), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[15]) );
  DFFR_X1 \program_cntr_out_reg[14]  ( .D(n566), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[14]) );
  DFFR_X1 \program_cntr_out_reg[13]  ( .D(n567), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[13]) );
  DFFR_X1 \program_cntr_out_reg[12]  ( .D(n568), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[12]) );
  DFFR_X1 \program_cntr_out_reg[11]  ( .D(n569), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[11]) );
  DFFR_X1 \program_cntr_out_reg[10]  ( .D(n570), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[10]) );
  DFFR_X1 \program_cntr_out_reg[9]  ( .D(n571), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[9]) );
  DFFR_X1 \program_cntr_out_reg[8]  ( .D(n572), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[8]) );
  DFFR_X1 \program_cntr_out_reg[7]  ( .D(n573), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[7]) );
  DFFR_X1 \program_cntr_out_reg[6]  ( .D(n574), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[6]) );
  DFFR_X1 \program_cntr_out_reg[5]  ( .D(n575), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[5]) );
  DFFR_X1 \program_cntr_out_reg[4]  ( .D(n576), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[4]) );
  DFFR_X1 \program_cntr_out_reg[3]  ( .D(n577), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[3]) );
  DFFR_X1 \program_cntr_out_reg[2]  ( .D(n578), .CK(clk_in), .RN(n143), .Q(
        program_cntr_out[2]) );
  DFFR_X1 \program_cntr_out_reg[1]  ( .D(n579), .CK(clk_in), .RN(n143), .Q(
        program_cntr_out[1]) );
  DFFR_X1 \program_cntr_out_reg[0]  ( .D(n580), .CK(clk_in), .RN(n143), .Q(
        program_cntr_out[0]) );
  DFFR_X1 \current_mask_out_reg[31]  ( .D(n581), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[31]) );
  DFFR_X1 \current_mask_out_reg[30]  ( .D(n582), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[30]) );
  DFFR_X1 \current_mask_out_reg[29]  ( .D(n583), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[29]) );
  DFFR_X1 \current_mask_out_reg[28]  ( .D(n584), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[28]) );
  DFFR_X1 \current_mask_out_reg[27]  ( .D(n585), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[27]) );
  DFFR_X1 \current_mask_out_reg[26]  ( .D(n586), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[26]) );
  DFFR_X1 \current_mask_out_reg[25]  ( .D(n587), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[25]) );
  DFFR_X1 \current_mask_out_reg[24]  ( .D(n588), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[24]) );
  DFFR_X1 \current_mask_out_reg[23]  ( .D(n589), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[23]) );
  DFFR_X1 \current_mask_out_reg[22]  ( .D(n590), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[22]) );
  DFFR_X1 \current_mask_out_reg[21]  ( .D(n591), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[21]) );
  DFFR_X1 \current_mask_out_reg[20]  ( .D(n592), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[20]) );
  DFFR_X1 \current_mask_out_reg[19]  ( .D(n593), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[19]) );
  DFFR_X1 \current_mask_out_reg[18]  ( .D(n594), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[18]) );
  DFFR_X1 \current_mask_out_reg[17]  ( .D(n595), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[17]) );
  DFFR_X1 \current_mask_out_reg[16]  ( .D(n596), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[16]) );
  DFFR_X1 \current_mask_out_reg[15]  ( .D(n597), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[15]) );
  DFFR_X1 \current_mask_out_reg[14]  ( .D(n598), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[14]) );
  DFFR_X1 \current_mask_out_reg[13]  ( .D(n599), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[13]) );
  DFFR_X1 \current_mask_out_reg[12]  ( .D(n600), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[12]) );
  DFFR_X1 \current_mask_out_reg[11]  ( .D(n601), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[11]) );
  DFFR_X1 \current_mask_out_reg[10]  ( .D(n602), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[10]) );
  DFFR_X1 \current_mask_out_reg[9]  ( .D(n603), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[9]) );
  DFFR_X1 \current_mask_out_reg[8]  ( .D(n604), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[8]) );
  DFFR_X1 \current_mask_out_reg[7]  ( .D(n605), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[7]) );
  DFFR_X1 \current_mask_out_reg[6]  ( .D(n606), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[6]) );
  DFFR_X1 \current_mask_out_reg[5]  ( .D(n607), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[5]) );
  DFFR_X1 \current_mask_out_reg[4]  ( .D(n608), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[4]) );
  DFFR_X1 \current_mask_out_reg[3]  ( .D(n609), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[3]) );
  DFFR_X1 \current_mask_out_reg[2]  ( .D(n610), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[2]) );
  DFFR_X1 \current_mask_out_reg[1]  ( .D(n611), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[1]) );
  DFFR_X1 \current_mask_out_reg[0]  ( .D(n612), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[0]) );
  DFFR_X1 \initial_mask_out_reg[31]  ( .D(n613), .CK(clk_in), .RN(n141), .Q(
        initial_mask_out[31]) );
  DFFR_X1 \initial_mask_out_reg[30]  ( .D(n614), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[30]) );
  DFFR_X1 \initial_mask_out_reg[29]  ( .D(n615), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[29]) );
  DFFR_X1 \initial_mask_out_reg[28]  ( .D(n616), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[28]) );
  DFFR_X1 \initial_mask_out_reg[27]  ( .D(n617), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[27]) );
  DFFR_X1 \initial_mask_out_reg[26]  ( .D(n618), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[26]) );
  DFFR_X1 \initial_mask_out_reg[25]  ( .D(n619), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[25]) );
  DFFR_X1 \initial_mask_out_reg[24]  ( .D(n620), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[24]) );
  DFFR_X1 \initial_mask_out_reg[23]  ( .D(n621), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[23]) );
  DFFR_X1 \initial_mask_out_reg[22]  ( .D(n622), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[22]) );
  DFFR_X1 \initial_mask_out_reg[21]  ( .D(n623), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[21]) );
  DFFR_X1 \initial_mask_out_reg[20]  ( .D(n624), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[20]) );
  DFFR_X1 \initial_mask_out_reg[19]  ( .D(n625), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[19]) );
  DFFR_X1 \initial_mask_out_reg[18]  ( .D(n626), .CK(clk_in), .RN(n139), .Q(
        initial_mask_out[18]) );
  DFFR_X1 \initial_mask_out_reg[17]  ( .D(n627), .CK(clk_in), .RN(n139), .Q(
        initial_mask_out[17]) );
  DFFR_X1 \initial_mask_out_reg[16]  ( .D(n628), .CK(clk_in), .RN(n139), .Q(
        initial_mask_out[16]) );
  DFFR_X1 \initial_mask_out_reg[15]  ( .D(n629), .CK(clk_in), .RN(n139), .Q(
        initial_mask_out[15]) );
  DFFR_X1 \initial_mask_out_reg[14]  ( .D(n630), .CK(clk_in), .RN(n139), .Q(
        initial_mask_out[14]) );
  DFFR_X1 \initial_mask_out_reg[13]  ( .D(n631), .CK(clk_in), .RN(n139), .Q(
        initial_mask_out[13]) );
  DFFR_X1 \warp_scheduler_next_state_reg[1]  ( .D(n422), .CK(clk_in), .RN(n139), .Q(warp_scheduler_next_state[1]), .QN(n182) );
  DFFR_X1 \warp_scheduler_state_machine_reg[1]  ( .D(n427), .CK(clk_in), .RN(
        n139), .Q(warp_scheduler_state_machine[1]), .QN(n166) );
  DFFR_X1 done_reg ( .D(n638), .CK(clk_in), .RN(n139), .Q(done) );
  DFFR_X1 \warp_state_wr_data_out_reg[0]  ( .D(n419), .CK(clk_in), .RN(n139), 
        .Q(warp_state_wr_data_out[0]) );
  DFFR_X1 warp_state_wr_en_out_reg ( .D(n420), .CK(clk_in), .RN(n139), .Q(
        warp_state_wr_en_out) );
  DFFR_X1 \warp_id_cnt_reg[1]  ( .D(n418), .CK(clk_in), .RN(n139), .Q(
        warp_id_cnt[1]), .QN(n179) );
  DFFR_X1 \warp_id_cnt_reg[4]  ( .D(n414), .CK(clk_in), .RN(n138), .Q(
        warp_id_cnt[4]), .QN(n170) );
  DFFR_X1 \warp_id_cnt_reg[3]  ( .D(n415), .CK(clk_in), .RN(n138), .Q(
        warp_id_cnt[3]), .QN(n177) );
  DFFR_X1 \warp_state_addr_out_reg[3]  ( .D(n405), .CK(clk_in), .RN(n138), .Q(
        warp_state_addr_out[3]) );
  DFFR_X1 \warp_pool_addr_out_reg[3]  ( .D(n410), .CK(clk_in), .RN(n138), .Q(
        warp_pool_addr_out[3]) );
  DFFR_X1 \warp_id_out_reg[3]  ( .D(n494), .CK(clk_in), .RN(n138), .Q(
        warp_id_out[3]) );
  DFFR_X1 \warp_id_cnt_reg[2]  ( .D(n416), .CK(clk_in), .RN(n138), .Q(
        warp_id_cnt[2]), .QN(n178) );
  DFFR_X1 \warp_state_addr_out_reg[2]  ( .D(n406), .CK(clk_in), .RN(n138), .Q(
        warp_state_addr_out[2]) );
  DFFR_X1 \warp_pool_addr_out_reg[2]  ( .D(n411), .CK(clk_in), .RN(n138), .Q(
        warp_pool_addr_out[2]) );
  DFFR_X1 \warp_id_out_reg[2]  ( .D(n495), .CK(clk_in), .RN(n138), .Q(
        warp_id_out[2]) );
  DFFR_X1 \warp_id_cnt_reg[0]  ( .D(n417), .CK(clk_in), .RN(n138), .Q(
        warp_id_cnt[0]), .QN(n180) );
  DFFR_X1 \warp_state_addr_out_reg[0]  ( .D(n408), .CK(clk_in), .RN(n138), .Q(
        warp_state_addr_out[0]) );
  DFFR_X1 \warp_pool_addr_out_reg[0]  ( .D(n413), .CK(clk_in), .RN(n138), .Q(
        warp_pool_addr_out[0]) );
  DFFR_X1 \warp_id_out_reg[0]  ( .D(n496), .CK(clk_in), .RN(n137), .Q(
        warp_id_out[0]) );
  DFFR_X1 \warp_state_addr_out_reg[4]  ( .D(n404), .CK(clk_in), .RN(n137), .Q(
        warp_state_addr_out[4]) );
  DFFR_X1 \warp_pool_addr_out_reg[4]  ( .D(n409), .CK(clk_in), .RN(n137), .Q(
        warp_pool_addr_out[4]) );
  DFFR_X1 \warp_id_out_reg[4]  ( .D(n493), .CK(clk_in), .RN(n137), .Q(
        warp_id_out[4]) );
  DFFR_X1 \warp_state_addr_out_reg[1]  ( .D(n407), .CK(clk_in), .RN(n137), .Q(
        warp_state_addr_out[1]) );
  DFFR_X1 \warp_pool_addr_out_reg[1]  ( .D(n412), .CK(clk_in), .RN(n137), .Q(
        warp_pool_addr_out[1]) );
  DFFR_X1 \warp_id_out_reg[1]  ( .D(n497), .CK(clk_in), .RN(n137), .Q(
        warp_id_out[1]) );
  DFFR_X1 pipeline_warpunit_done_reg ( .D(n426), .CK(clk_in), .RN(n137), .Q(
        pipeline_warpunit_done) );
  DFFR_X1 fetch_en_reg ( .D(n424), .CK(clk_in), .RN(n137), .Q(fetch_en) );
  DFFR_X1 \warp_lane_cnt_reg[0]  ( .D(n423), .CK(clk_in), .RN(n137), .Q(
        warp_lane_cnt[0]), .QN(n169) );
  DFFR_X1 \warp_lane_id_out_reg[0]  ( .D(n498), .CK(clk_in), .RN(n137), .Q(
        warp_lane_id_out[0]) );
  DFFR_X1 \warp_lane_id_out_reg[1]  ( .D(n499), .CK(clk_in), .RN(n137), .Q(
        warp_lane_id_out[1]) );
  NAND2_X1 U382 ( .A1(warp_state_addr_out[4]), .A2(n632), .ZN(n190) );
  NAND2_X1 U383 ( .A1(warp_state_addr_out[3]), .A2(n632), .ZN(n192) );
  NAND2_X1 U384 ( .A1(warp_state_addr_out[2]), .A2(n632), .ZN(n194) );
  NAND2_X1 U385 ( .A1(warp_state_addr_out[1]), .A2(n632), .ZN(n196) );
  NAND2_X1 U386 ( .A1(warp_state_addr_out[0]), .A2(n632), .ZN(n198) );
  NAND2_X1 U387 ( .A1(n202), .A2(n203), .ZN(n199) );
  NAND2_X1 U388 ( .A1(warp_pool_addr_out[4]), .A2(n202), .ZN(n204) );
  NAND2_X1 U389 ( .A1(N73), .A2(n205), .ZN(n189) );
  NAND2_X1 U390 ( .A1(warp_pool_addr_out[3]), .A2(n202), .ZN(n206) );
  NAND2_X1 U391 ( .A1(N72), .A2(n205), .ZN(n191) );
  NAND2_X1 U392 ( .A1(warp_pool_addr_out[2]), .A2(n202), .ZN(n207) );
  NAND2_X1 U393 ( .A1(N71), .A2(n205), .ZN(n193) );
  NAND2_X1 U394 ( .A1(warp_pool_addr_out[1]), .A2(n202), .ZN(n208) );
  NAND2_X1 U395 ( .A1(N70), .A2(n205), .ZN(n195) );
  NAND2_X1 U396 ( .A1(warp_pool_addr_out[0]), .A2(n202), .ZN(n209) );
  NAND2_X1 U397 ( .A1(n180), .A2(n205), .ZN(n197) );
  NAND2_X1 U398 ( .A1(n210), .A2(n221), .ZN(n213) );
  NAND3_X1 U399 ( .A1(n222), .A2(n492), .A3(n223), .ZN(n221) );
  NAND2_X1 U400 ( .A1(n225), .A2(n226), .ZN(n210) );
  NAND2_X1 U401 ( .A1(warp_state_wr_data_out[0]), .A2(n131), .ZN(n228) );
  NAND2_X1 U402 ( .A1(warp_state_wr_en_out), .A2(n229), .ZN(n230) );
  NAND3_X1 U403 ( .A1(n237), .A2(n169), .A3(n239), .ZN(n238) );
  NAND2_X1 U404 ( .A1(fetch_en), .A2(n240), .ZN(n242) );
  NAND3_X1 U405 ( .A1(n239), .A2(n237), .A3(n248), .ZN(n247) );
  NAND2_X1 U406 ( .A1(pipeline_warpunit_done), .A2(n387), .ZN(n388) );
  NAND3_X1 U407 ( .A1(n166), .A2(n161), .A3(n167), .ZN(n392) );
  NAND2_X1 U408 ( .A1(n640), .A2(n231), .ZN(n201) );
  NAND3_X1 U409 ( .A1(warp_scheduler_state_machine[1]), .A2(n167), .A3(
        warp_scheduler_state_machine[2]), .ZN(n231) );
  NAND3_X1 U410 ( .A1(n220), .A2(n232), .A3(n226), .ZN(n235) );
  NAND2_X1 U411 ( .A1(n449), .A2(n403), .ZN(n232) );
  NAND2_X1 U414 ( .A1(n252), .A2(n200), .ZN(n203) );
  warps_done_lut uWarpsDoneLUT ( .clk_in(clk_in), .host_reset(host_reset), 
        .num_warps_in(num_warps_in), .warps_done_mask(warps_done_mask) );
  warp_scheduler_SHMEM_ADDR_SIZE14_DW01_cmp6_1 eq_164 ( .A(warps_done_mask_in), 
        .B(warps_done_mask), .TC(1'b0), .EQ(N52) );
  HA_X1 \r149/U1_1_1  ( .A(warp_id_cnt[1]), .B(warp_id_cnt[0]), .CO(
        \r149/carry[2] ), .S(N70) );
  HA_X1 \r149/U1_1_2  ( .A(warp_id_cnt[2]), .B(\r149/carry[2] ), .CO(
        \r149/carry[3] ), .S(N71) );
  HA_X1 \r149/U1_1_3  ( .A(warp_id_cnt[3]), .B(\r149/carry[3] ), .CO(
        \r149/carry[4] ), .S(N72) );
  NOR3_X1 U133 ( .A1(n167), .A2(warp_scheduler_state_machine[2]), .A3(n166), 
        .ZN(n200) );
  NOR3_X1 U134 ( .A1(warp_scheduler_state_machine[0]), .A2(
        warp_scheduler_state_machine[2]), .A3(n166), .ZN(n244) );
  NOR3_X1 U135 ( .A1(warp_scheduler_state_machine[0]), .A2(
        warp_scheduler_state_machine[1]), .A3(n161), .ZN(n220) );
  AND2_X1 U136 ( .A1(n250), .A2(n203), .ZN(n130) );
  INV_X1 U137 ( .A(n448), .ZN(n154) );
  INV_X1 U138 ( .A(n449), .ZN(n156) );
  INV_X1 U139 ( .A(n447), .ZN(n152) );
  INV_X1 U140 ( .A(n449), .ZN(n157) );
  BUF_X1 U141 ( .A(n450), .Z(n448) );
  BUF_X1 U142 ( .A(n450), .Z(n449) );
  BUF_X1 U143 ( .A(n450), .Z(n447) );
  BUF_X1 U144 ( .A(n451), .Z(n446) );
  BUF_X1 U145 ( .A(n451), .Z(n445) );
  BUF_X1 U146 ( .A(n451), .Z(n444) );
  BUF_X1 U147 ( .A(n452), .Z(n443) );
  BUF_X1 U148 ( .A(n452), .Z(n442) );
  BUF_X1 U149 ( .A(n452), .Z(n441) );
  BUF_X1 U150 ( .A(n453), .Z(n440) );
  BUF_X1 U151 ( .A(n453), .Z(n439) );
  BUF_X1 U152 ( .A(n453), .Z(n438) );
  BUF_X1 U153 ( .A(n454), .Z(n437) );
  BUF_X1 U154 ( .A(n454), .Z(n436) );
  BUF_X1 U155 ( .A(n454), .Z(n435) );
  BUF_X1 U156 ( .A(n455), .Z(n434) );
  BUF_X1 U157 ( .A(n455), .Z(n433) );
  BUF_X1 U158 ( .A(n455), .Z(n432) );
  BUF_X1 U159 ( .A(n456), .Z(n212) );
  BUF_X1 U160 ( .A(n456), .Z(n187) );
  BUF_X1 U161 ( .A(n457), .Z(n186) );
  BUF_X1 U162 ( .A(n457), .Z(n185) );
  BUF_X1 U163 ( .A(n457), .Z(n184) );
  BUF_X1 U164 ( .A(n458), .Z(n176) );
  BUF_X1 U165 ( .A(n458), .Z(n175) );
  BUF_X1 U166 ( .A(n458), .Z(n174) );
  BUF_X1 U167 ( .A(n459), .Z(n173) );
  BUF_X1 U168 ( .A(n459), .Z(n172) );
  BUF_X1 U169 ( .A(n456), .Z(n431) );
  BUF_X1 U170 ( .A(n459), .Z(n171) );
  BUF_X1 U171 ( .A(n460), .Z(n165) );
  BUF_X1 U172 ( .A(n460), .Z(n164) );
  BUF_X1 U173 ( .A(n460), .Z(n163) );
  BUF_X1 U174 ( .A(n461), .Z(n162) );
  BUF_X1 U175 ( .A(n461), .Z(n160) );
  BUF_X1 U176 ( .A(n461), .Z(n159) );
  BUF_X1 U177 ( .A(n462), .Z(n158) );
  BUF_X1 U178 ( .A(n453), .Z(n462) );
  BUF_X1 U179 ( .A(n455), .Z(n457) );
  BUF_X1 U180 ( .A(n453), .Z(n458) );
  BUF_X1 U181 ( .A(n452), .Z(n456) );
  BUF_X1 U182 ( .A(n454), .Z(n459) );
  BUF_X1 U183 ( .A(n453), .Z(n460) );
  BUF_X1 U184 ( .A(n454), .Z(n461) );
  BUF_X1 U185 ( .A(n130), .Z(n450) );
  BUF_X1 U186 ( .A(n130), .Z(n451) );
  BUF_X1 U187 ( .A(n130), .Z(n452) );
  BUF_X1 U188 ( .A(n130), .Z(n453) );
  BUF_X1 U189 ( .A(n130), .Z(n454) );
  BUF_X1 U190 ( .A(n130), .Z(n455) );
  INV_X1 U191 ( .A(n199), .ZN(n632) );
  INV_X1 U192 ( .A(N52), .ZN(n492) );
  NOR2_X1 U193 ( .A1(n492), .A2(n635), .ZN(n397) );
  INV_X1 U194 ( .A(n478), .ZN(n486) );
  AND2_X1 U195 ( .A1(n639), .A2(n210), .ZN(n202) );
  INV_X1 U196 ( .A(n201), .ZN(n639) );
  NOR2_X1 U197 ( .A1(n635), .A2(n648), .ZN(n243) );
  NOR2_X1 U198 ( .A1(n642), .A2(n641), .ZN(n205) );
  AND3_X1 U199 ( .A1(n640), .A2(n203), .A3(n641), .ZN(n131) );
  INV_X1 U200 ( .A(n227), .ZN(n636) );
  INV_X1 U201 ( .A(n223), .ZN(n633) );
  BUF_X1 U202 ( .A(n132), .Z(n134) );
  BUF_X1 U203 ( .A(n132), .Z(n135) );
  BUF_X1 U204 ( .A(n132), .Z(n136) );
  OAI211_X1 U205 ( .C1(n219), .C2(n220), .A(n213), .B(N67), .ZN(n214) );
  INV_X1 U206 ( .A(n220), .ZN(n641) );
  NOR2_X1 U207 ( .A1(n244), .A2(n225), .ZN(n250) );
  INV_X1 U208 ( .A(n398), .ZN(n490) );
  INV_X1 U209 ( .A(n232), .ZN(n491) );
  INV_X1 U210 ( .A(N67), .ZN(n642) );
  INV_X1 U211 ( .A(N66), .ZN(n484) );
  OAI21_X1 U212 ( .B1(n200), .B2(n201), .A(n199), .ZN(n188) );
  OAI21_X1 U213 ( .B1(n249), .B2(n635), .A(n250), .ZN(n237) );
  NOR2_X1 U214 ( .A1(n251), .A2(n252), .ZN(n249) );
  NOR3_X1 U215 ( .A1(n253), .A2(N52), .A3(n254), .ZN(n251) );
  NOR2_X1 U216 ( .A1(n641), .A2(n226), .ZN(n234) );
  NOR2_X1 U217 ( .A1(n244), .A2(n200), .ZN(n227) );
  NOR2_X1 U218 ( .A1(n635), .A2(n254), .ZN(n223) );
  NOR2_X1 U219 ( .A1(n220), .A2(n243), .ZN(n390) );
  NOR2_X1 U220 ( .A1(n647), .A2(n649), .ZN(n253) );
  INV_X1 U221 ( .A(n200), .ZN(n635) );
  INV_X1 U222 ( .A(n244), .ZN(n640) );
  NAND4_X1 U223 ( .A1(n391), .A2(n637), .A3(n640), .A4(n392), .ZN(n245) );
  OR3_X1 U224 ( .A1(n253), .A2(N52), .A3(n635), .ZN(n391) );
  INV_X1 U225 ( .A(n393), .ZN(n637) );
  OR3_X1 U226 ( .A1(n243), .A2(n234), .A3(n244), .ZN(n239) );
  INV_X1 U227 ( .A(n468), .ZN(n485) );
  INV_X1 U228 ( .A(n254), .ZN(n648) );
  NOR2_X1 U229 ( .A1(host_reset), .A2(reset), .ZN(n132) );
  OAI22_X1 U230 ( .A1(warp_state_rd_data_in[1]), .A2(N94), .B1(
        pipeline_stall_in), .B2(n224), .ZN(n222) );
  INV_X1 U231 ( .A(n477), .ZN(n488) );
  NAND4_X1 U232 ( .A1(warp_state_rd_data_in[1]), .A2(n200), .A3(n492), .A4(
        n647), .ZN(n403) );
  OAI211_X1 U233 ( .C1(pipeline_stall_in), .C2(n390), .A(n639), .B(n402), .ZN(
        n398) );
  AOI221_X1 U234 ( .B1(n223), .B2(n649), .C1(warp_scheduler_state_machine[0]), 
        .C2(n166), .A(n397), .ZN(n402) );
  INV_X1 U235 ( .A(n332), .ZN(n577) );
  AOI22_X1 U236 ( .A1(program_cntr_out[3]), .A2(n432), .B1(N418), .B2(n154), 
        .ZN(n332) );
  NOR3_X1 U237 ( .A1(N52), .A2(pipeline_stall_in), .A3(n648), .ZN(n252) );
  NOR2_X1 U238 ( .A1(n641), .A2(pipeline_stall_in), .ZN(n225) );
  XOR2_X1 U239 ( .A(num_warps_in[3]), .B(n465), .Z(n133) );
  OAI221_X1 U240 ( .B1(n491), .B2(n633), .C1(n232), .C2(n182), .A(n235), .ZN(
        n422) );
  OAI22_X1 U241 ( .A1(n180), .A2(n213), .B1(warp_id_cnt[0]), .B2(n214), .ZN(
        n417) );
  OAI22_X1 U242 ( .A1(n178), .A2(n213), .B1(n645), .B2(n214), .ZN(n416) );
  INV_X1 U243 ( .A(N71), .ZN(n645) );
  OAI22_X1 U244 ( .A1(n177), .A2(n213), .B1(n644), .B2(n214), .ZN(n415) );
  INV_X1 U245 ( .A(N72), .ZN(n644) );
  OAI22_X1 U246 ( .A1(n170), .A2(n213), .B1(n643), .B2(n214), .ZN(n414) );
  INV_X1 U247 ( .A(N73), .ZN(n643) );
  OAI22_X1 U248 ( .A1(n179), .A2(n213), .B1(n646), .B2(n214), .ZN(n418) );
  INV_X1 U249 ( .A(N70), .ZN(n646) );
  OAI22_X1 U250 ( .A1(n232), .A2(n181), .B1(n491), .B2(n233), .ZN(n421) );
  NOR2_X1 U251 ( .A1(n234), .A2(n636), .ZN(n233) );
  INV_X1 U252 ( .A(n481), .ZN(n487) );
  AOI21_X1 U253 ( .B1(warp_state_rd_data_in[1]), .B2(n642), .A(n219), .ZN(n224) );
  INV_X1 U254 ( .A(n474), .ZN(n489) );
  OAI21_X1 U255 ( .B1(n232), .B2(n183), .A(n235), .ZN(n430) );
  INV_X1 U256 ( .A(num_warps_in[2]), .ZN(n467) );
  NAND4_X1 U257 ( .A1(n633), .A2(n392), .A3(n231), .A4(n396), .ZN(n427) );
  AOI221_X1 U258 ( .B1(n490), .B2(warp_scheduler_state_machine[1]), .C1(n393), 
        .C2(warp_scheduler_next_state[1]), .A(n397), .ZN(n396) );
  INV_X1 U259 ( .A(n335), .ZN(n580) );
  AOI22_X1 U260 ( .A1(program_cntr_out[0]), .A2(n433), .B1(N415), .B2(n154), 
        .ZN(n335) );
  INV_X1 U261 ( .A(n334), .ZN(n579) );
  AOI22_X1 U262 ( .A1(program_cntr_out[1]), .A2(n432), .B1(N416), .B2(n156), 
        .ZN(n334) );
  INV_X1 U263 ( .A(n333), .ZN(n578) );
  AOI22_X1 U264 ( .A1(program_cntr_out[2]), .A2(n432), .B1(N417), .B2(n151), 
        .ZN(n333) );
  INV_X1 U265 ( .A(n331), .ZN(n576) );
  AOI22_X1 U266 ( .A1(program_cntr_out[4]), .A2(n432), .B1(N419), .B2(n154), 
        .ZN(n331) );
  INV_X1 U267 ( .A(n330), .ZN(n575) );
  AOI22_X1 U268 ( .A1(program_cntr_out[5]), .A2(n431), .B1(N420), .B2(n154), 
        .ZN(n330) );
  INV_X1 U269 ( .A(n329), .ZN(n574) );
  AOI22_X1 U270 ( .A1(program_cntr_out[6]), .A2(n431), .B1(N421), .B2(n154), 
        .ZN(n329) );
  INV_X1 U271 ( .A(n328), .ZN(n573) );
  AOI22_X1 U272 ( .A1(program_cntr_out[7]), .A2(n431), .B1(N422), .B2(n154), 
        .ZN(n328) );
  INV_X1 U273 ( .A(n327), .ZN(n572) );
  AOI22_X1 U274 ( .A1(program_cntr_out[8]), .A2(n212), .B1(N423), .B2(n154), 
        .ZN(n327) );
  INV_X1 U275 ( .A(n326), .ZN(n571) );
  AOI22_X1 U276 ( .A1(program_cntr_out[9]), .A2(n212), .B1(N424), .B2(n154), 
        .ZN(n326) );
  INV_X1 U277 ( .A(n325), .ZN(n570) );
  AOI22_X1 U278 ( .A1(program_cntr_out[10]), .A2(n212), .B1(N425), .B2(n154), 
        .ZN(n325) );
  INV_X1 U279 ( .A(n324), .ZN(n569) );
  AOI22_X1 U280 ( .A1(program_cntr_out[11]), .A2(n212), .B1(N426), .B2(n154), 
        .ZN(n324) );
  INV_X1 U281 ( .A(n323), .ZN(n568) );
  AOI22_X1 U282 ( .A1(program_cntr_out[12]), .A2(n187), .B1(N427), .B2(n155), 
        .ZN(n323) );
  INV_X1 U283 ( .A(n322), .ZN(n567) );
  AOI22_X1 U284 ( .A1(program_cntr_out[13]), .A2(n187), .B1(N428), .B2(n155), 
        .ZN(n322) );
  INV_X1 U285 ( .A(n321), .ZN(n566) );
  AOI22_X1 U286 ( .A1(program_cntr_out[14]), .A2(n187), .B1(N429), .B2(n155), 
        .ZN(n321) );
  INV_X1 U287 ( .A(n320), .ZN(n565) );
  AOI22_X1 U288 ( .A1(program_cntr_out[15]), .A2(n187), .B1(N430), .B2(n155), 
        .ZN(n320) );
  INV_X1 U289 ( .A(n319), .ZN(n564) );
  AOI22_X1 U290 ( .A1(program_cntr_out[16]), .A2(n186), .B1(N431), .B2(n155), 
        .ZN(n319) );
  INV_X1 U291 ( .A(n318), .ZN(n563) );
  AOI22_X1 U292 ( .A1(program_cntr_out[17]), .A2(n186), .B1(N432), .B2(n155), 
        .ZN(n318) );
  INV_X1 U293 ( .A(n377), .ZN(n622) );
  AOI22_X1 U294 ( .A1(initial_mask_out[22]), .A2(n443), .B1(N372), .B2(n151), 
        .ZN(n377) );
  INV_X1 U295 ( .A(n376), .ZN(n621) );
  AOI22_X1 U296 ( .A1(initial_mask_out[23]), .A2(n443), .B1(N373), .B2(n151), 
        .ZN(n376) );
  INV_X1 U297 ( .A(n375), .ZN(n620) );
  AOI22_X1 U298 ( .A1(initial_mask_out[24]), .A2(n443), .B1(N375), .B2(n151), 
        .ZN(n375) );
  INV_X1 U299 ( .A(n374), .ZN(n619) );
  AOI22_X1 U300 ( .A1(initial_mask_out[25]), .A2(n442), .B1(N376), .B2(n151), 
        .ZN(n374) );
  INV_X1 U301 ( .A(n373), .ZN(n618) );
  AOI22_X1 U302 ( .A1(initial_mask_out[26]), .A2(n442), .B1(N377), .B2(n151), 
        .ZN(n373) );
  INV_X1 U303 ( .A(n372), .ZN(n617) );
  AOI22_X1 U304 ( .A1(initial_mask_out[27]), .A2(n442), .B1(N378), .B2(n151), 
        .ZN(n372) );
  INV_X1 U305 ( .A(n371), .ZN(n616) );
  AOI22_X1 U306 ( .A1(initial_mask_out[28]), .A2(n442), .B1(N379), .B2(n151), 
        .ZN(n371) );
  INV_X1 U307 ( .A(n370), .ZN(n615) );
  AOI22_X1 U308 ( .A1(initial_mask_out[29]), .A2(n441), .B1(N380), .B2(n151), 
        .ZN(n370) );
  INV_X1 U309 ( .A(n369), .ZN(n614) );
  AOI22_X1 U310 ( .A1(initial_mask_out[30]), .A2(n441), .B1(N381), .B2(n151), 
        .ZN(n369) );
  INV_X1 U311 ( .A(n350), .ZN(n595) );
  AOI22_X1 U312 ( .A1(current_mask_out[17]), .A2(n436), .B1(N400), .B2(n153), 
        .ZN(n350) );
  INV_X1 U313 ( .A(n349), .ZN(n594) );
  AOI22_X1 U314 ( .A1(current_mask_out[18]), .A2(n436), .B1(N401), .B2(n153), 
        .ZN(n349) );
  INV_X1 U315 ( .A(n348), .ZN(n593) );
  AOI22_X1 U316 ( .A1(current_mask_out[19]), .A2(n436), .B1(N402), .B2(n153), 
        .ZN(n348) );
  INV_X1 U317 ( .A(n347), .ZN(n592) );
  AOI22_X1 U318 ( .A1(current_mask_out[20]), .A2(n436), .B1(N403), .B2(n153), 
        .ZN(n347) );
  INV_X1 U319 ( .A(n346), .ZN(n591) );
  AOI22_X1 U320 ( .A1(current_mask_out[21]), .A2(n435), .B1(N404), .B2(n153), 
        .ZN(n346) );
  INV_X1 U321 ( .A(n345), .ZN(n590) );
  AOI22_X1 U322 ( .A1(current_mask_out[22]), .A2(n435), .B1(N405), .B2(n153), 
        .ZN(n345) );
  INV_X1 U323 ( .A(n344), .ZN(n589) );
  AOI22_X1 U324 ( .A1(current_mask_out[23]), .A2(n435), .B1(N406), .B2(n153), 
        .ZN(n344) );
  INV_X1 U325 ( .A(n343), .ZN(n588) );
  AOI22_X1 U326 ( .A1(current_mask_out[24]), .A2(n435), .B1(N407), .B2(n153), 
        .ZN(n343) );
  INV_X1 U327 ( .A(n342), .ZN(n587) );
  AOI22_X1 U328 ( .A1(current_mask_out[25]), .A2(n434), .B1(N408), .B2(n153), 
        .ZN(n342) );
  INV_X1 U329 ( .A(n341), .ZN(n586) );
  AOI22_X1 U330 ( .A1(current_mask_out[26]), .A2(n434), .B1(N409), .B2(n151), 
        .ZN(n341) );
  INV_X1 U331 ( .A(n340), .ZN(n585) );
  AOI22_X1 U332 ( .A1(current_mask_out[27]), .A2(n434), .B1(N410), .B2(n154), 
        .ZN(n340) );
  INV_X1 U333 ( .A(n339), .ZN(n584) );
  AOI22_X1 U334 ( .A1(current_mask_out[28]), .A2(n434), .B1(N411), .B2(n154), 
        .ZN(n339) );
  INV_X1 U335 ( .A(n338), .ZN(n583) );
  AOI22_X1 U336 ( .A1(current_mask_out[29]), .A2(n433), .B1(N412), .B2(n151), 
        .ZN(n338) );
  INV_X1 U337 ( .A(n337), .ZN(n582) );
  AOI22_X1 U338 ( .A1(current_mask_out[30]), .A2(n433), .B1(N413), .B2(n153), 
        .ZN(n337) );
  INV_X1 U339 ( .A(n336), .ZN(n581) );
  AOI22_X1 U340 ( .A1(current_mask_out[31]), .A2(n433), .B1(N414), .B2(n151), 
        .ZN(n336) );
  INV_X1 U341 ( .A(n317), .ZN(n562) );
  AOI22_X1 U342 ( .A1(program_cntr_out[18]), .A2(n186), .B1(N433), .B2(n155), 
        .ZN(n317) );
  INV_X1 U343 ( .A(n316), .ZN(n561) );
  AOI22_X1 U344 ( .A1(program_cntr_out[19]), .A2(n186), .B1(N434), .B2(n155), 
        .ZN(n316) );
  INV_X1 U345 ( .A(n315), .ZN(n560) );
  AOI22_X1 U346 ( .A1(program_cntr_out[20]), .A2(n185), .B1(N435), .B2(n155), 
        .ZN(n315) );
  INV_X1 U347 ( .A(n314), .ZN(n559) );
  AOI22_X1 U348 ( .A1(program_cntr_out[21]), .A2(n185), .B1(N436), .B2(n156), 
        .ZN(n314) );
  INV_X1 U349 ( .A(n313), .ZN(n558) );
  AOI22_X1 U350 ( .A1(program_cntr_out[22]), .A2(n185), .B1(N437), .B2(n156), 
        .ZN(n313) );
  INV_X1 U351 ( .A(n312), .ZN(n557) );
  AOI22_X1 U352 ( .A1(program_cntr_out[23]), .A2(n185), .B1(N438), .B2(n156), 
        .ZN(n312) );
  INV_X1 U353 ( .A(n311), .ZN(n556) );
  AOI22_X1 U354 ( .A1(program_cntr_out[24]), .A2(n184), .B1(N439), .B2(n156), 
        .ZN(n311) );
  INV_X1 U355 ( .A(n310), .ZN(n555) );
  AOI22_X1 U356 ( .A1(program_cntr_out[25]), .A2(n184), .B1(N440), .B2(n156), 
        .ZN(n310) );
  INV_X1 U357 ( .A(n309), .ZN(n554) );
  AOI22_X1 U358 ( .A1(program_cntr_out[26]), .A2(n184), .B1(N441), .B2(n156), 
        .ZN(n309) );
  INV_X1 U359 ( .A(n308), .ZN(n553) );
  AOI22_X1 U360 ( .A1(program_cntr_out[27]), .A2(n184), .B1(N442), .B2(n156), 
        .ZN(n308) );
  INV_X1 U361 ( .A(n307), .ZN(n552) );
  AOI22_X1 U362 ( .A1(program_cntr_out[28]), .A2(n176), .B1(N443), .B2(n156), 
        .ZN(n307) );
  INV_X1 U363 ( .A(n306), .ZN(n551) );
  AOI22_X1 U364 ( .A1(program_cntr_out[29]), .A2(n176), .B1(N444), .B2(n156), 
        .ZN(n306) );
  INV_X1 U365 ( .A(n305), .ZN(n550) );
  AOI22_X1 U366 ( .A1(program_cntr_out[30]), .A2(n176), .B1(N445), .B2(n151), 
        .ZN(n305) );
  INV_X1 U367 ( .A(n246), .ZN(n499) );
  AOI22_X1 U368 ( .A1(n157), .A2(warp_lane_cnt[1]), .B1(n446), .B2(
        warp_lane_id_out[1]), .ZN(n246) );
  INV_X1 U369 ( .A(n236), .ZN(n498) );
  AOI22_X1 U370 ( .A1(n157), .A2(warp_lane_cnt[0]), .B1(n446), .B2(
        warp_lane_id_out[0]), .ZN(n236) );
  INV_X1 U371 ( .A(n218), .ZN(n497) );
  AOI22_X1 U372 ( .A1(n157), .A2(warp_id_cnt[1]), .B1(n446), .B2(
        warp_id_out[1]), .ZN(n218) );
  INV_X1 U373 ( .A(n304), .ZN(n549) );
  AOI22_X1 U374 ( .A1(program_cntr_out[31]), .A2(n176), .B1(N446), .B2(n154), 
        .ZN(n304) );
  INV_X1 U375 ( .A(n211), .ZN(n493) );
  AOI22_X1 U376 ( .A1(n152), .A2(warp_id_cnt[4]), .B1(n447), .B2(
        warp_id_out[4]), .ZN(n211) );
  INV_X1 U377 ( .A(n217), .ZN(n496) );
  AOI22_X1 U378 ( .A1(n157), .A2(warp_id_cnt[0]), .B1(n447), .B2(
        warp_id_out[0]), .ZN(n217) );
  INV_X1 U379 ( .A(n216), .ZN(n495) );
  AOI22_X1 U380 ( .A1(n152), .A2(warp_id_cnt[2]), .B1(n446), .B2(
        warp_id_out[2]), .ZN(n216) );
  INV_X1 U381 ( .A(n215), .ZN(n494) );
  AOI22_X1 U412 ( .A1(n157), .A2(warp_id_cnt[3]), .B1(n447), .B2(
        warp_id_out[3]), .ZN(n215) );
  INV_X1 U413 ( .A(n303), .ZN(n548) );
  AOI22_X1 U415 ( .A1(gprs_size_out[0]), .A2(n175), .B1(N447), .B2(n153), .ZN(
        n303) );
  INV_X1 U416 ( .A(n302), .ZN(n547) );
  AOI22_X1 U417 ( .A1(gprs_size_out[1]), .A2(n175), .B1(N448), .B2(n154), .ZN(
        n302) );
  INV_X1 U418 ( .A(n301), .ZN(n546) );
  AOI22_X1 U419 ( .A1(gprs_size_out[2]), .A2(n175), .B1(N449), .B2(n151), .ZN(
        n301) );
  INV_X1 U420 ( .A(n300), .ZN(n545) );
  AOI22_X1 U421 ( .A1(gprs_size_out[3]), .A2(n175), .B1(N450), .B2(n151), .ZN(
        n300) );
  INV_X1 U422 ( .A(n299), .ZN(n544) );
  AOI22_X1 U423 ( .A1(gprs_size_out[4]), .A2(n174), .B1(N451), .B2(n153), .ZN(
        n299) );
  INV_X1 U424 ( .A(n298), .ZN(n543) );
  AOI22_X1 U425 ( .A1(gprs_size_out[5]), .A2(n174), .B1(N452), .B2(n154), .ZN(
        n298) );
  INV_X1 U426 ( .A(n297), .ZN(n542) );
  AOI22_X1 U427 ( .A1(gprs_size_out[6]), .A2(n174), .B1(N453), .B2(n151), .ZN(
        n297) );
  INV_X1 U428 ( .A(n296), .ZN(n541) );
  AOI22_X1 U429 ( .A1(gprs_size_out[7]), .A2(n174), .B1(N454), .B2(n155), .ZN(
        n296) );
  INV_X1 U430 ( .A(n295), .ZN(n540) );
  AOI22_X1 U431 ( .A1(gprs_size_out[8]), .A2(n173), .B1(N455), .B2(n157), .ZN(
        n295) );
  INV_X1 U432 ( .A(n294), .ZN(n539) );
  AOI22_X1 U433 ( .A1(shmem_base_addr_out[0]), .A2(n173), .B1(N321), .B2(n156), 
        .ZN(n294) );
  INV_X1 U434 ( .A(n293), .ZN(n538) );
  AOI22_X1 U435 ( .A1(shmem_base_addr_out[1]), .A2(n173), .B1(N322), .B2(n152), 
        .ZN(n293) );
  INV_X1 U436 ( .A(n292), .ZN(n537) );
  AOI22_X1 U437 ( .A1(shmem_base_addr_out[2]), .A2(n173), .B1(N323), .B2(n153), 
        .ZN(n292) );
  INV_X1 U438 ( .A(n291), .ZN(n536) );
  AOI22_X1 U439 ( .A1(shmem_base_addr_out[3]), .A2(n172), .B1(N324), .B2(n153), 
        .ZN(n291) );
  INV_X1 U440 ( .A(n290), .ZN(n535) );
  AOI22_X1 U441 ( .A1(shmem_base_addr_out[4]), .A2(n172), .B1(N325), .B2(n155), 
        .ZN(n290) );
  INV_X1 U442 ( .A(n289), .ZN(n534) );
  AOI22_X1 U443 ( .A1(shmem_base_addr_out[5]), .A2(n172), .B1(N326), .B2(n157), 
        .ZN(n289) );
  INV_X1 U444 ( .A(n288), .ZN(n533) );
  AOI22_X1 U445 ( .A1(shmem_base_addr_out[6]), .A2(n172), .B1(N327), .B2(n156), 
        .ZN(n288) );
  INV_X1 U446 ( .A(n287), .ZN(n532) );
  AOI22_X1 U447 ( .A1(shmem_base_addr_out[7]), .A2(n171), .B1(N328), .B2(n151), 
        .ZN(n287) );
  INV_X1 U448 ( .A(n286), .ZN(n531) );
  AOI22_X1 U449 ( .A1(shmem_base_addr_out[8]), .A2(n171), .B1(N329), .B2(n152), 
        .ZN(n286) );
  INV_X1 U450 ( .A(n285), .ZN(n530) );
  AOI22_X1 U451 ( .A1(shmem_base_addr_out[9]), .A2(n431), .B1(N330), .B2(n153), 
        .ZN(n285) );
  INV_X1 U452 ( .A(n284), .ZN(n529) );
  AOI22_X1 U453 ( .A1(shmem_base_addr_out[10]), .A2(n171), .B1(N331), .B2(n154), .ZN(n284) );
  INV_X1 U454 ( .A(n283), .ZN(n528) );
  AOI22_X1 U455 ( .A1(shmem_base_addr_out[11]), .A2(n171), .B1(N332), .B2(n151), .ZN(n283) );
  INV_X1 U456 ( .A(n282), .ZN(n527) );
  AOI22_X1 U457 ( .A1(shmem_base_addr_out[12]), .A2(n165), .B1(N333), .B2(n152), .ZN(n282) );
  INV_X1 U458 ( .A(n281), .ZN(n526) );
  AOI22_X1 U459 ( .A1(shmem_base_addr_out[13]), .A2(n165), .B1(N334), .B2(n155), .ZN(n281) );
  INV_X1 U460 ( .A(n280), .ZN(n525) );
  AOI22_X1 U461 ( .A1(cta_id_out[0]), .A2(n165), .B1(N335), .B2(n156), .ZN(
        n280) );
  INV_X1 U462 ( .A(n279), .ZN(n524) );
  AOI22_X1 U463 ( .A1(cta_id_out[1]), .A2(n165), .B1(N336), .B2(n157), .ZN(
        n279) );
  INV_X1 U464 ( .A(n278), .ZN(n523) );
  AOI22_X1 U465 ( .A1(cta_id_out[2]), .A2(n164), .B1(N337), .B2(n151), .ZN(
        n278) );
  INV_X1 U466 ( .A(n277), .ZN(n522) );
  AOI22_X1 U467 ( .A1(cta_id_out[3]), .A2(n164), .B1(N338), .B2(n153), .ZN(
        n277) );
  INV_X1 U468 ( .A(n276), .ZN(n521) );
  AOI22_X1 U469 ( .A1(gprs_base_addr_out[0]), .A2(n164), .B1(N339), .B2(n153), 
        .ZN(n276) );
  INV_X1 U470 ( .A(n275), .ZN(n520) );
  AOI22_X1 U471 ( .A1(gprs_base_addr_out[1]), .A2(n164), .B1(N340), .B2(n151), 
        .ZN(n275) );
  INV_X1 U472 ( .A(n274), .ZN(n519) );
  AOI22_X1 U473 ( .A1(gprs_base_addr_out[2]), .A2(n163), .B1(N341), .B2(n154), 
        .ZN(n274) );
  INV_X1 U474 ( .A(n273), .ZN(n518) );
  AOI22_X1 U475 ( .A1(gprs_base_addr_out[3]), .A2(n163), .B1(N342), .B2(n154), 
        .ZN(n273) );
  INV_X1 U476 ( .A(n272), .ZN(n517) );
  AOI22_X1 U477 ( .A1(gprs_base_addr_out[4]), .A2(n163), .B1(N343), .B2(n154), 
        .ZN(n272) );
  INV_X1 U478 ( .A(n271), .ZN(n516) );
  AOI22_X1 U479 ( .A1(gprs_base_addr_out[5]), .A2(n163), .B1(N344), .B2(n154), 
        .ZN(n271) );
  INV_X1 U480 ( .A(n270), .ZN(n515) );
  AOI22_X1 U481 ( .A1(gprs_base_addr_out[6]), .A2(n162), .B1(N345), .B2(n153), 
        .ZN(n270) );
  INV_X1 U482 ( .A(n269), .ZN(n514) );
  AOI22_X1 U483 ( .A1(gprs_base_addr_out[7]), .A2(n162), .B1(N346), .B2(n155), 
        .ZN(n269) );
  INV_X1 U484 ( .A(n268), .ZN(n513) );
  AOI22_X1 U485 ( .A1(gprs_base_addr_out[8]), .A2(n162), .B1(N347), .B2(n155), 
        .ZN(n268) );
  INV_X1 U486 ( .A(n267), .ZN(n512) );
  AOI22_X1 U487 ( .A1(initial_mask_out[0]), .A2(n162), .B1(N348), .B2(n153), 
        .ZN(n267) );
  INV_X1 U488 ( .A(n266), .ZN(n511) );
  AOI22_X1 U489 ( .A1(initial_mask_out[1]), .A2(n160), .B1(N349), .B2(n153), 
        .ZN(n266) );
  INV_X1 U490 ( .A(n265), .ZN(n510) );
  AOI22_X1 U491 ( .A1(initial_mask_out[2]), .A2(n160), .B1(N350), .B2(n157), 
        .ZN(n265) );
  INV_X1 U492 ( .A(n264), .ZN(n509) );
  AOI22_X1 U493 ( .A1(initial_mask_out[3]), .A2(n160), .B1(N351), .B2(n156), 
        .ZN(n264) );
  INV_X1 U494 ( .A(n263), .ZN(n508) );
  AOI22_X1 U495 ( .A1(initial_mask_out[4]), .A2(n160), .B1(N352), .B2(n157), 
        .ZN(n263) );
  INV_X1 U496 ( .A(n262), .ZN(n507) );
  AOI22_X1 U497 ( .A1(initial_mask_out[5]), .A2(n159), .B1(N353), .B2(n155), 
        .ZN(n262) );
  INV_X1 U498 ( .A(n261), .ZN(n506) );
  AOI22_X1 U499 ( .A1(initial_mask_out[6]), .A2(n159), .B1(N354), .B2(n154), 
        .ZN(n261) );
  INV_X1 U500 ( .A(n386), .ZN(n631) );
  AOI22_X1 U501 ( .A1(initial_mask_out[13]), .A2(n445), .B1(N362), .B2(n156), 
        .ZN(n386) );
  INV_X1 U502 ( .A(n385), .ZN(n630) );
  AOI22_X1 U503 ( .A1(initial_mask_out[14]), .A2(n445), .B1(N364), .B2(n155), 
        .ZN(n385) );
  INV_X1 U504 ( .A(n384), .ZN(n629) );
  AOI22_X1 U505 ( .A1(initial_mask_out[15]), .A2(n445), .B1(N365), .B2(n153), 
        .ZN(n384) );
  INV_X1 U506 ( .A(n383), .ZN(n628) );
  AOI22_X1 U507 ( .A1(initial_mask_out[16]), .A2(n445), .B1(N366), .B2(n157), 
        .ZN(n383) );
  INV_X1 U508 ( .A(n382), .ZN(n627) );
  AOI22_X1 U509 ( .A1(initial_mask_out[17]), .A2(n444), .B1(N367), .B2(n152), 
        .ZN(n382) );
  INV_X1 U510 ( .A(n381), .ZN(n626) );
  AOI22_X1 U511 ( .A1(initial_mask_out[18]), .A2(n444), .B1(N368), .B2(n155), 
        .ZN(n381) );
  INV_X1 U512 ( .A(n380), .ZN(n625) );
  AOI22_X1 U513 ( .A1(initial_mask_out[19]), .A2(n444), .B1(N369), .B2(n156), 
        .ZN(n380) );
  INV_X1 U514 ( .A(n379), .ZN(n624) );
  AOI22_X1 U515 ( .A1(initial_mask_out[20]), .A2(n444), .B1(N370), .B2(n157), 
        .ZN(n379) );
  INV_X1 U516 ( .A(n378), .ZN(n623) );
  AOI22_X1 U517 ( .A1(initial_mask_out[21]), .A2(n443), .B1(N371), .B2(n157), 
        .ZN(n378) );
  INV_X1 U518 ( .A(n368), .ZN(n613) );
  AOI22_X1 U519 ( .A1(initial_mask_out[31]), .A2(n441), .B1(N382), .B2(n152), 
        .ZN(n368) );
  INV_X1 U520 ( .A(n367), .ZN(n612) );
  AOI22_X1 U521 ( .A1(current_mask_out[0]), .A2(n441), .B1(N383), .B2(n152), 
        .ZN(n367) );
  INV_X1 U522 ( .A(n366), .ZN(n611) );
  AOI22_X1 U523 ( .A1(current_mask_out[1]), .A2(n440), .B1(N384), .B2(n152), 
        .ZN(n366) );
  INV_X1 U524 ( .A(n365), .ZN(n610) );
  AOI22_X1 U525 ( .A1(current_mask_out[2]), .A2(n440), .B1(N385), .B2(n152), 
        .ZN(n365) );
  INV_X1 U526 ( .A(n364), .ZN(n609) );
  AOI22_X1 U527 ( .A1(current_mask_out[3]), .A2(n440), .B1(N386), .B2(n152), 
        .ZN(n364) );
  INV_X1 U528 ( .A(n363), .ZN(n608) );
  AOI22_X1 U529 ( .A1(current_mask_out[4]), .A2(n440), .B1(N387), .B2(n152), 
        .ZN(n363) );
  INV_X1 U530 ( .A(n362), .ZN(n607) );
  AOI22_X1 U531 ( .A1(current_mask_out[5]), .A2(n439), .B1(N388), .B2(n152), 
        .ZN(n362) );
  INV_X1 U532 ( .A(n361), .ZN(n606) );
  AOI22_X1 U533 ( .A1(current_mask_out[6]), .A2(n439), .B1(N389), .B2(n152), 
        .ZN(n361) );
  INV_X1 U534 ( .A(n360), .ZN(n605) );
  AOI22_X1 U535 ( .A1(current_mask_out[7]), .A2(n439), .B1(N390), .B2(n152), 
        .ZN(n360) );
  INV_X1 U536 ( .A(n359), .ZN(n604) );
  AOI22_X1 U537 ( .A1(current_mask_out[8]), .A2(n439), .B1(N391), .B2(n152), 
        .ZN(n359) );
  INV_X1 U538 ( .A(n358), .ZN(n603) );
  AOI22_X1 U539 ( .A1(current_mask_out[9]), .A2(n438), .B1(N392), .B2(n152), 
        .ZN(n358) );
  INV_X1 U540 ( .A(n357), .ZN(n602) );
  AOI22_X1 U541 ( .A1(current_mask_out[10]), .A2(n438), .B1(N393), .B2(n152), 
        .ZN(n357) );
  INV_X1 U542 ( .A(n356), .ZN(n601) );
  AOI22_X1 U543 ( .A1(current_mask_out[11]), .A2(n438), .B1(N394), .B2(n155), 
        .ZN(n356) );
  INV_X1 U544 ( .A(n355), .ZN(n600) );
  AOI22_X1 U545 ( .A1(current_mask_out[12]), .A2(n438), .B1(N395), .B2(n152), 
        .ZN(n355) );
  INV_X1 U546 ( .A(n354), .ZN(n599) );
  AOI22_X1 U547 ( .A1(current_mask_out[13]), .A2(n437), .B1(N396), .B2(n156), 
        .ZN(n354) );
  INV_X1 U548 ( .A(n353), .ZN(n598) );
  AOI22_X1 U549 ( .A1(current_mask_out[14]), .A2(n437), .B1(N397), .B2(n156), 
        .ZN(n353) );
  INV_X1 U550 ( .A(n352), .ZN(n597) );
  AOI22_X1 U551 ( .A1(current_mask_out[15]), .A2(n437), .B1(N398), .B2(n156), 
        .ZN(n352) );
  INV_X1 U552 ( .A(n351), .ZN(n596) );
  AOI22_X1 U553 ( .A1(current_mask_out[16]), .A2(n437), .B1(N399), .B2(n155), 
        .ZN(n351) );
  INV_X1 U554 ( .A(n260), .ZN(n505) );
  AOI22_X1 U555 ( .A1(initial_mask_out[7]), .A2(n159), .B1(N355), .B2(n157), 
        .ZN(n260) );
  INV_X1 U556 ( .A(n259), .ZN(n504) );
  AOI22_X1 U557 ( .A1(initial_mask_out[8]), .A2(n159), .B1(N356), .B2(n157), 
        .ZN(n259) );
  INV_X1 U558 ( .A(n258), .ZN(n503) );
  AOI22_X1 U559 ( .A1(initial_mask_out[9]), .A2(n158), .B1(N357), .B2(n157), 
        .ZN(n258) );
  INV_X1 U560 ( .A(n257), .ZN(n502) );
  AOI22_X1 U561 ( .A1(initial_mask_out[10]), .A2(n158), .B1(N358), .B2(n157), 
        .ZN(n257) );
  INV_X1 U562 ( .A(n256), .ZN(n501) );
  AOI22_X1 U563 ( .A1(initial_mask_out[11]), .A2(n158), .B1(N359), .B2(n157), 
        .ZN(n256) );
  INV_X1 U564 ( .A(n255), .ZN(n500) );
  AOI22_X1 U565 ( .A1(initial_mask_out[12]), .A2(n158), .B1(N360), .B2(n157), 
        .ZN(n255) );
  NOR3_X1 U566 ( .A1(n167), .A2(warp_scheduler_state_machine[1]), .A3(n161), 
        .ZN(n393) );
  OAI221_X1 U567 ( .B1(n188), .B2(n179), .C1(n632), .C2(n195), .A(n196), .ZN(
        n407) );
  OAI221_X1 U568 ( .B1(n188), .B2(n170), .C1(n632), .C2(n189), .A(n190), .ZN(
        n404) );
  OAI221_X1 U569 ( .B1(n188), .B2(n180), .C1(n632), .C2(n197), .A(n198), .ZN(
        n408) );
  OAI221_X1 U570 ( .B1(n188), .B2(n178), .C1(n632), .C2(n193), .A(n194), .ZN(
        n406) );
  OAI221_X1 U571 ( .B1(n188), .B2(n177), .C1(n632), .C2(n191), .A(n192), .ZN(
        n405) );
  OAI221_X1 U572 ( .B1(n639), .B2(n179), .C1(n202), .C2(n195), .A(n208), .ZN(
        n412) );
  OAI221_X1 U573 ( .B1(n639), .B2(n170), .C1(n202), .C2(n189), .A(n204), .ZN(
        n409) );
  OAI221_X1 U574 ( .B1(n639), .B2(n180), .C1(n202), .C2(n197), .A(n209), .ZN(
        n413) );
  OAI221_X1 U575 ( .B1(n639), .B2(n178), .C1(n202), .C2(n193), .A(n207), .ZN(
        n411) );
  OAI221_X1 U576 ( .B1(n639), .B2(n177), .C1(n202), .C2(n191), .A(n206), .ZN(
        n410) );
  NOR2_X1 U577 ( .A1(n168), .A2(n169), .ZN(n226) );
  OAI22_X1 U578 ( .A1(n161), .A2(n398), .B1(n490), .B2(n401), .ZN(n429) );
  AOI211_X1 U579 ( .C1(n393), .C2(warp_scheduler_next_state[2]), .A(n636), .B(
        n220), .ZN(n401) );
  OAI22_X1 U580 ( .A1(n167), .A2(n398), .B1(n490), .B2(n399), .ZN(n428) );
  AND3_X1 U581 ( .A1(n400), .A2(n639), .A3(n390), .ZN(n399) );
  AOI21_X1 U582 ( .B1(n393), .B2(warp_scheduler_next_state[0]), .A(n397), .ZN(
        n400) );
  OAI21_X1 U583 ( .B1(n390), .B2(pipeline_stall_in), .A(n640), .ZN(n389) );
  INV_X1 U584 ( .A(pipeline_stall_in), .ZN(n647) );
  OAI21_X1 U585 ( .B1(n227), .B2(n229), .A(n230), .ZN(n420) );
  AND3_X1 U586 ( .A1(n231), .A2(n131), .A3(n637), .ZN(n229) );
  OAI21_X1 U587 ( .B1(n131), .B2(n227), .A(n228), .ZN(n419) );
  OAI21_X1 U588 ( .B1(n387), .B2(n634), .A(n388), .ZN(n426) );
  INV_X1 U589 ( .A(n389), .ZN(n634) );
  NOR2_X1 U590 ( .A1(n245), .A2(n220), .ZN(n387) );
  OAI21_X1 U591 ( .B1(n240), .B2(n241), .A(n242), .ZN(n424) );
  AOI21_X1 U592 ( .B1(n243), .B2(n647), .A(n244), .ZN(n241) );
  NOR3_X1 U593 ( .A1(n225), .A2(n234), .A3(n245), .ZN(n240) );
  OAI21_X1 U594 ( .B1(n168), .B2(n237), .A(n247), .ZN(n425) );
  XNOR2_X1 U595 ( .A(n168), .B(warp_lane_cnt[0]), .ZN(n248) );
  OAI21_X1 U596 ( .B1(n169), .B2(n237), .A(n238), .ZN(n423) );
  INV_X1 U597 ( .A(n394), .ZN(n638) );
  AOI21_X1 U598 ( .B1(n392), .B2(done), .A(n395), .ZN(n394) );
  NOR3_X1 U599 ( .A1(n166), .A2(n167), .A3(n161), .ZN(n395) );
  NOR2_X1 U600 ( .A1(warp_state_rd_data_in[1]), .A2(warp_state_rd_data_in[0]), 
        .ZN(n254) );
  AND2_X1 U601 ( .A1(warp_state_rd_data_in[0]), .A2(warp_state_rd_data_in[1]), 
        .ZN(n219) );
  INV_X1 U602 ( .A(warp_state_rd_data_in[1]), .ZN(n649) );
  CLKBUF_X1 U603 ( .A(n134), .Z(n137) );
  CLKBUF_X1 U604 ( .A(n134), .Z(n138) );
  CLKBUF_X1 U605 ( .A(n134), .Z(n139) );
  CLKBUF_X1 U606 ( .A(n134), .Z(n140) );
  CLKBUF_X1 U607 ( .A(n134), .Z(n141) );
  CLKBUF_X1 U608 ( .A(n134), .Z(n142) );
  CLKBUF_X1 U609 ( .A(n135), .Z(n143) );
  CLKBUF_X1 U610 ( .A(n135), .Z(n144) );
  CLKBUF_X1 U611 ( .A(n135), .Z(n145) );
  CLKBUF_X1 U612 ( .A(n135), .Z(n146) );
  CLKBUF_X1 U613 ( .A(n135), .Z(n147) );
  CLKBUF_X1 U614 ( .A(n135), .Z(n148) );
  CLKBUF_X1 U615 ( .A(n136), .Z(n149) );
  CLKBUF_X1 U616 ( .A(n136), .Z(n150) );
  INV_X1 U617 ( .A(n448), .ZN(n151) );
  INV_X1 U618 ( .A(n448), .ZN(n153) );
  INV_X1 U619 ( .A(n449), .ZN(n155) );
  NOR2_X1 U620 ( .A1(num_warps_in[1]), .A2(num_warps_in[0]), .ZN(n464) );
  AOI21_X1 U621 ( .B1(num_warps_in[0]), .B2(num_warps_in[1]), .A(n464), .ZN(
        n463) );
  INV_X1 U622 ( .A(n463), .ZN(N63) );
  NAND2_X1 U623 ( .A1(n464), .A2(n467), .ZN(n465) );
  OAI21_X1 U624 ( .B1(n464), .B2(n467), .A(n465), .ZN(N64) );
  NOR2_X1 U625 ( .A1(num_warps_in[3]), .A2(n465), .ZN(n466) );
  XOR2_X1 U626 ( .A(num_warps_in[4]), .B(n466), .Z(N66) );
  XOR2_X1 U627 ( .A(\r149/carry[4] ), .B(warp_id_cnt[4]), .Z(N73) );
  NOR2_X1 U628 ( .A1(n178), .A2(N64), .ZN(n469) );
  NAND2_X1 U629 ( .A1(warp_id_cnt[3]), .A2(n133), .ZN(n481) );
  NOR2_X1 U630 ( .A1(n469), .A2(n487), .ZN(n472) );
  NAND2_X1 U631 ( .A1(warp_id_cnt[0]), .A2(num_warps_in[0]), .ZN(n468) );
  OAI21_X1 U632 ( .B1(n179), .B2(n468), .A(N63), .ZN(n470) );
  NAND2_X1 U633 ( .A1(N64), .A2(n178), .ZN(n478) );
  NOR2_X1 U634 ( .A1(n469), .A2(n486), .ZN(n475) );
  OAI211_X1 U635 ( .C1(warp_id_cnt[1]), .C2(n485), .A(n470), .B(n475), .ZN(
        n471) );
  NOR2_X1 U636 ( .A1(n133), .A2(warp_id_cnt[3]), .ZN(n477) );
  AOI21_X1 U637 ( .B1(n472), .B2(n471), .A(n477), .ZN(n473) );
  XNOR2_X1 U638 ( .A(warp_id_cnt[4]), .B(N66), .ZN(n480) );
  AOI22_X1 U639 ( .A1(n473), .A2(n480), .B1(warp_id_cnt[4]), .B2(n484), .ZN(
        N94) );
  NOR2_X1 U640 ( .A1(num_warps_in[0]), .A2(warp_id_cnt[0]), .ZN(n476) );
  AOI21_X1 U641 ( .B1(n179), .B2(n476), .A(N63), .ZN(n474) );
  OAI211_X1 U642 ( .C1(n476), .C2(n179), .A(n489), .B(n475), .ZN(n479) );
  NAND3_X1 U643 ( .A1(n479), .A2(n478), .A3(n488), .ZN(n482) );
  NAND3_X1 U644 ( .A1(n482), .A2(n481), .A3(n480), .ZN(n483) );
  OAI21_X1 U645 ( .B1(warp_id_cnt[4]), .B2(n484), .A(n483), .ZN(N67) );
endmodule




module warp_unit ( clk_in, host_reset, warp_scheduler_reset, 
        warp_generator_en, pipeline_write_done, pipeline_stall_in, 
        threads_per_block_in, num_blocks_in, warps_per_block_in, 
        shared_mem_base_addr_in, shared_mem_size_in, gprs_size_in, block_x_in, 
        block_y_in, block_z_in, grid_x_in, grid_y_in, block_idx_in, warp_id_in, 
        warp_lane_id_in, cta_id_in, initial_mask_in, current_mask_in, 
        shmem_base_addr_in, gprs_base_addr_in, next_pc_in, warp_state_in, 
        program_cntr_out, warp_id_out, warp_lane_id_out, cta_id_out, 
        initial_mask_out, current_mask_out, shmem_base_addr_out, gprs_size_out, 
        gprs_base_addr_out, num_warps_out, warp_generator_done, 
        pipeline_stall_out, warp_scheduler_done, pipeline_warpunit_done, 
        fetch_en );
  input [11:0] threads_per_block_in;
  input [3:0] num_blocks_in;
  input [5:0] warps_per_block_in;
  input [31:0] shared_mem_base_addr_in;
  input [31:0] shared_mem_size_in;
  input [8:0] gprs_size_in;
  input [15:0] block_x_in;
  input [15:0] block_y_in;
  input [15:0] block_z_in;
  input [15:0] grid_x_in;
  input [15:0] grid_y_in;
  input [15:0] block_idx_in;
  input [4:0] warp_id_in;
  input [1:0] warp_lane_id_in;
  input [3:0] cta_id_in;
  input [31:0] initial_mask_in;
  input [31:0] current_mask_in;
  input [13:0] shmem_base_addr_in;
  input [8:0] gprs_base_addr_in;
  input [31:0] next_pc_in;
  input [1:0] warp_state_in;
  output [31:0] program_cntr_out;
  output [4:0] warp_id_out;
  output [1:0] warp_lane_id_out;
  output [3:0] cta_id_out;
  output [31:0] initial_mask_out;
  output [31:0] current_mask_out;
  output [13:0] shmem_base_addr_out;
  output [8:0] gprs_size_out;
  output [8:0] gprs_base_addr_out;
  output [4:0] num_warps_out;
  input clk_in, host_reset, warp_scheduler_reset, warp_generator_en,
         pipeline_write_done, pipeline_stall_in;
  output warp_generator_done, pipeline_stall_out, warp_scheduler_done,
         pipeline_warpunit_done, fetch_en;
  wire   warp_gen_pool_wr_en, warp_gen_state_wr_en,
         \warp_gen_fence_regs_wr_cta_id[31><3] ,
         \warp_gen_fence_regs_wr_cta_id[31><2] ,
         \warp_gen_fence_regs_wr_cta_id[31><1] ,
         \warp_gen_fence_regs_wr_cta_id[31><0] ,
         \warp_gen_fence_regs_wr_cta_id[30><3] ,
         \warp_gen_fence_regs_wr_cta_id[30><2] ,
         \warp_gen_fence_regs_wr_cta_id[30><1] ,
         \warp_gen_fence_regs_wr_cta_id[30><0] ,
         \warp_gen_fence_regs_wr_cta_id[29><3] ,
         \warp_gen_fence_regs_wr_cta_id[29><2] ,
         \warp_gen_fence_regs_wr_cta_id[29><1] ,
         \warp_gen_fence_regs_wr_cta_id[29><0] ,
         \warp_gen_fence_regs_wr_cta_id[28><3] ,
         \warp_gen_fence_regs_wr_cta_id[28><2] ,
         \warp_gen_fence_regs_wr_cta_id[28><1] ,
         \warp_gen_fence_regs_wr_cta_id[28><0] ,
         \warp_gen_fence_regs_wr_cta_id[27><3] ,
         \warp_gen_fence_regs_wr_cta_id[27><2] ,
         \warp_gen_fence_regs_wr_cta_id[27><1] ,
         \warp_gen_fence_regs_wr_cta_id[27><0] ,
         \warp_gen_fence_regs_wr_cta_id[26><3] ,
         \warp_gen_fence_regs_wr_cta_id[26><2] ,
         \warp_gen_fence_regs_wr_cta_id[26><1] ,
         \warp_gen_fence_regs_wr_cta_id[26><0] ,
         \warp_gen_fence_regs_wr_cta_id[25><3] ,
         \warp_gen_fence_regs_wr_cta_id[25><2] ,
         \warp_gen_fence_regs_wr_cta_id[25><1] ,
         \warp_gen_fence_regs_wr_cta_id[25><0] ,
         \warp_gen_fence_regs_wr_cta_id[24><3] ,
         \warp_gen_fence_regs_wr_cta_id[24><2] ,
         \warp_gen_fence_regs_wr_cta_id[24><1] ,
         \warp_gen_fence_regs_wr_cta_id[24><0] ,
         \warp_gen_fence_regs_wr_cta_id[23><3] ,
         \warp_gen_fence_regs_wr_cta_id[23><2] ,
         \warp_gen_fence_regs_wr_cta_id[23><1] ,
         \warp_gen_fence_regs_wr_cta_id[23><0] ,
         \warp_gen_fence_regs_wr_cta_id[22><3] ,
         \warp_gen_fence_regs_wr_cta_id[22><2] ,
         \warp_gen_fence_regs_wr_cta_id[22><1] ,
         \warp_gen_fence_regs_wr_cta_id[22><0] ,
         \warp_gen_fence_regs_wr_cta_id[21><3] ,
         \warp_gen_fence_regs_wr_cta_id[21><2] ,
         \warp_gen_fence_regs_wr_cta_id[21><1] ,
         \warp_gen_fence_regs_wr_cta_id[21><0] ,
         \warp_gen_fence_regs_wr_cta_id[20><3] ,
         \warp_gen_fence_regs_wr_cta_id[20><2] ,
         \warp_gen_fence_regs_wr_cta_id[20><1] ,
         \warp_gen_fence_regs_wr_cta_id[20><0] ,
         \warp_gen_fence_regs_wr_cta_id[19><3] ,
         \warp_gen_fence_regs_wr_cta_id[19><2] ,
         \warp_gen_fence_regs_wr_cta_id[19><1] ,
         \warp_gen_fence_regs_wr_cta_id[19><0] ,
         \warp_gen_fence_regs_wr_cta_id[18><3] ,
         \warp_gen_fence_regs_wr_cta_id[18><2] ,
         \warp_gen_fence_regs_wr_cta_id[18><1] ,
         \warp_gen_fence_regs_wr_cta_id[18><0] ,
         \warp_gen_fence_regs_wr_cta_id[17><3] ,
         \warp_gen_fence_regs_wr_cta_id[17><2] ,
         \warp_gen_fence_regs_wr_cta_id[17><1] ,
         \warp_gen_fence_regs_wr_cta_id[17><0] ,
         \warp_gen_fence_regs_wr_cta_id[16><3] ,
         \warp_gen_fence_regs_wr_cta_id[16><2] ,
         \warp_gen_fence_regs_wr_cta_id[16><1] ,
         \warp_gen_fence_regs_wr_cta_id[16><0] ,
         \warp_gen_fence_regs_wr_cta_id[15><3] ,
         \warp_gen_fence_regs_wr_cta_id[15><2] ,
         \warp_gen_fence_regs_wr_cta_id[15><1] ,
         \warp_gen_fence_regs_wr_cta_id[15><0] ,
         \warp_gen_fence_regs_wr_cta_id[14><3] ,
         \warp_gen_fence_regs_wr_cta_id[14><2] ,
         \warp_gen_fence_regs_wr_cta_id[14><1] ,
         \warp_gen_fence_regs_wr_cta_id[14><0] ,
         \warp_gen_fence_regs_wr_cta_id[13><3] ,
         \warp_gen_fence_regs_wr_cta_id[13><2] ,
         \warp_gen_fence_regs_wr_cta_id[13><1] ,
         \warp_gen_fence_regs_wr_cta_id[13><0] ,
         \warp_gen_fence_regs_wr_cta_id[12><3] ,
         \warp_gen_fence_regs_wr_cta_id[12><2] ,
         \warp_gen_fence_regs_wr_cta_id[12><1] ,
         \warp_gen_fence_regs_wr_cta_id[12><0] ,
         \warp_gen_fence_regs_wr_cta_id[11><3] ,
         \warp_gen_fence_regs_wr_cta_id[11><2] ,
         \warp_gen_fence_regs_wr_cta_id[11><1] ,
         \warp_gen_fence_regs_wr_cta_id[11><0] ,
         \warp_gen_fence_regs_wr_cta_id[10><3] ,
         \warp_gen_fence_regs_wr_cta_id[10><2] ,
         \warp_gen_fence_regs_wr_cta_id[10><1] ,
         \warp_gen_fence_regs_wr_cta_id[10><0] ,
         \warp_gen_fence_regs_wr_cta_id[9><3] ,
         \warp_gen_fence_regs_wr_cta_id[9><2] ,
         \warp_gen_fence_regs_wr_cta_id[9><1] ,
         \warp_gen_fence_regs_wr_cta_id[9><0] ,
         \warp_gen_fence_regs_wr_cta_id[8><3] ,
         \warp_gen_fence_regs_wr_cta_id[8><2] ,
         \warp_gen_fence_regs_wr_cta_id[8><1] ,
         \warp_gen_fence_regs_wr_cta_id[8><0] ,
         \warp_gen_fence_regs_wr_cta_id[7><3] ,
         \warp_gen_fence_regs_wr_cta_id[7><2] ,
         \warp_gen_fence_regs_wr_cta_id[7><1] ,
         \warp_gen_fence_regs_wr_cta_id[7><0] ,
         \warp_gen_fence_regs_wr_cta_id[6><3] ,
         \warp_gen_fence_regs_wr_cta_id[6><2] ,
         \warp_gen_fence_regs_wr_cta_id[6><1] ,
         \warp_gen_fence_regs_wr_cta_id[6><0] ,
         \warp_gen_fence_regs_wr_cta_id[5><3] ,
         \warp_gen_fence_regs_wr_cta_id[5><2] ,
         \warp_gen_fence_regs_wr_cta_id[5><1] ,
         \warp_gen_fence_regs_wr_cta_id[5><0] ,
         \warp_gen_fence_regs_wr_cta_id[4><3] ,
         \warp_gen_fence_regs_wr_cta_id[4><2] ,
         \warp_gen_fence_regs_wr_cta_id[4><1] ,
         \warp_gen_fence_regs_wr_cta_id[4><0] ,
         \warp_gen_fence_regs_wr_cta_id[3><3] ,
         \warp_gen_fence_regs_wr_cta_id[3><2] ,
         \warp_gen_fence_regs_wr_cta_id[3><1] ,
         \warp_gen_fence_regs_wr_cta_id[3><0] ,
         \warp_gen_fence_regs_wr_cta_id[2><3] ,
         \warp_gen_fence_regs_wr_cta_id[2><2] ,
         \warp_gen_fence_regs_wr_cta_id[2><1] ,
         \warp_gen_fence_regs_wr_cta_id[2><0] ,
         \warp_gen_fence_regs_wr_cta_id[1><3] ,
         \warp_gen_fence_regs_wr_cta_id[1><2] ,
         \warp_gen_fence_regs_wr_cta_id[1><1] ,
         \warp_gen_fence_regs_wr_cta_id[1><0] ,
         \warp_gen_fence_regs_wr_cta_id[0><3] ,
         \warp_gen_fence_regs_wr_cta_id[0><2] ,
         \warp_gen_fence_regs_wr_cta_id[0><1] ,
         \warp_gen_fence_regs_wr_cta_id[0><0] , warp_sched_state_wr_en,
         \warp_sched_state_wr_data[0] , warp_pool_wr_en_b, warp_state_wr_en_b,
         \warp_checker_fence_regs_rd_cta_id[31><3] ,
         \warp_checker_fence_regs_rd_cta_id[31><2] ,
         \warp_checker_fence_regs_rd_cta_id[31><1] ,
         \warp_checker_fence_regs_rd_cta_id[31><0] ,
         \warp_checker_fence_regs_rd_cta_id[30><3] ,
         \warp_checker_fence_regs_rd_cta_id[30><2] ,
         \warp_checker_fence_regs_rd_cta_id[30><1] ,
         \warp_checker_fence_regs_rd_cta_id[30><0] ,
         \warp_checker_fence_regs_rd_cta_id[29><3] ,
         \warp_checker_fence_regs_rd_cta_id[29><2] ,
         \warp_checker_fence_regs_rd_cta_id[29><1] ,
         \warp_checker_fence_regs_rd_cta_id[29><0] ,
         \warp_checker_fence_regs_rd_cta_id[28><3] ,
         \warp_checker_fence_regs_rd_cta_id[28><2] ,
         \warp_checker_fence_regs_rd_cta_id[28><1] ,
         \warp_checker_fence_regs_rd_cta_id[28><0] ,
         \warp_checker_fence_regs_rd_cta_id[27><3] ,
         \warp_checker_fence_regs_rd_cta_id[27><2] ,
         \warp_checker_fence_regs_rd_cta_id[27><1] ,
         \warp_checker_fence_regs_rd_cta_id[27><0] ,
         \warp_checker_fence_regs_rd_cta_id[26><3] ,
         \warp_checker_fence_regs_rd_cta_id[26><2] ,
         \warp_checker_fence_regs_rd_cta_id[26><1] ,
         \warp_checker_fence_regs_rd_cta_id[26><0] ,
         \warp_checker_fence_regs_rd_cta_id[25><3] ,
         \warp_checker_fence_regs_rd_cta_id[25><2] ,
         \warp_checker_fence_regs_rd_cta_id[25><1] ,
         \warp_checker_fence_regs_rd_cta_id[25><0] ,
         \warp_checker_fence_regs_rd_cta_id[24><3] ,
         \warp_checker_fence_regs_rd_cta_id[24><2] ,
         \warp_checker_fence_regs_rd_cta_id[24><1] ,
         \warp_checker_fence_regs_rd_cta_id[24><0] ,
         \warp_checker_fence_regs_rd_cta_id[23><3] ,
         \warp_checker_fence_regs_rd_cta_id[23><2] ,
         \warp_checker_fence_regs_rd_cta_id[23><1] ,
         \warp_checker_fence_regs_rd_cta_id[23><0] ,
         \warp_checker_fence_regs_rd_cta_id[22><3] ,
         \warp_checker_fence_regs_rd_cta_id[22><2] ,
         \warp_checker_fence_regs_rd_cta_id[22><1] ,
         \warp_checker_fence_regs_rd_cta_id[22><0] ,
         \warp_checker_fence_regs_rd_cta_id[21><3] ,
         \warp_checker_fence_regs_rd_cta_id[21><2] ,
         \warp_checker_fence_regs_rd_cta_id[21><1] ,
         \warp_checker_fence_regs_rd_cta_id[21><0] ,
         \warp_checker_fence_regs_rd_cta_id[20><3] ,
         \warp_checker_fence_regs_rd_cta_id[20><2] ,
         \warp_checker_fence_regs_rd_cta_id[20><1] ,
         \warp_checker_fence_regs_rd_cta_id[20><0] ,
         \warp_checker_fence_regs_rd_cta_id[19><3] ,
         \warp_checker_fence_regs_rd_cta_id[19><2] ,
         \warp_checker_fence_regs_rd_cta_id[19><1] ,
         \warp_checker_fence_regs_rd_cta_id[19><0] ,
         \warp_checker_fence_regs_rd_cta_id[18><3] ,
         \warp_checker_fence_regs_rd_cta_id[18><2] ,
         \warp_checker_fence_regs_rd_cta_id[18><1] ,
         \warp_checker_fence_regs_rd_cta_id[18><0] ,
         \warp_checker_fence_regs_rd_cta_id[17><3] ,
         \warp_checker_fence_regs_rd_cta_id[17><2] ,
         \warp_checker_fence_regs_rd_cta_id[17><1] ,
         \warp_checker_fence_regs_rd_cta_id[17><0] ,
         \warp_checker_fence_regs_rd_cta_id[16><3] ,
         \warp_checker_fence_regs_rd_cta_id[16><2] ,
         \warp_checker_fence_regs_rd_cta_id[16><1] ,
         \warp_checker_fence_regs_rd_cta_id[16><0] ,
         \warp_checker_fence_regs_rd_cta_id[15><3] ,
         \warp_checker_fence_regs_rd_cta_id[15><2] ,
         \warp_checker_fence_regs_rd_cta_id[15><1] ,
         \warp_checker_fence_regs_rd_cta_id[15><0] ,
         \warp_checker_fence_regs_rd_cta_id[14><3] ,
         \warp_checker_fence_regs_rd_cta_id[14><2] ,
         \warp_checker_fence_regs_rd_cta_id[14><1] ,
         \warp_checker_fence_regs_rd_cta_id[14><0] ,
         \warp_checker_fence_regs_rd_cta_id[13><3] ,
         \warp_checker_fence_regs_rd_cta_id[13><2] ,
         \warp_checker_fence_regs_rd_cta_id[13><1] ,
         \warp_checker_fence_regs_rd_cta_id[13><0] ,
         \warp_checker_fence_regs_rd_cta_id[12><3] ,
         \warp_checker_fence_regs_rd_cta_id[12><2] ,
         \warp_checker_fence_regs_rd_cta_id[12><1] ,
         \warp_checker_fence_regs_rd_cta_id[12><0] ,
         \warp_checker_fence_regs_rd_cta_id[11><3] ,
         \warp_checker_fence_regs_rd_cta_id[11><2] ,
         \warp_checker_fence_regs_rd_cta_id[11><1] ,
         \warp_checker_fence_regs_rd_cta_id[11><0] ,
         \warp_checker_fence_regs_rd_cta_id[10><3] ,
         \warp_checker_fence_regs_rd_cta_id[10><2] ,
         \warp_checker_fence_regs_rd_cta_id[10><1] ,
         \warp_checker_fence_regs_rd_cta_id[10><0] ,
         \warp_checker_fence_regs_rd_cta_id[9><3] ,
         \warp_checker_fence_regs_rd_cta_id[9><2] ,
         \warp_checker_fence_regs_rd_cta_id[9><1] ,
         \warp_checker_fence_regs_rd_cta_id[9><0] ,
         \warp_checker_fence_regs_rd_cta_id[8><3] ,
         \warp_checker_fence_regs_rd_cta_id[8><2] ,
         \warp_checker_fence_regs_rd_cta_id[8><1] ,
         \warp_checker_fence_regs_rd_cta_id[8><0] ,
         \warp_checker_fence_regs_rd_cta_id[7><3] ,
         \warp_checker_fence_regs_rd_cta_id[7><2] ,
         \warp_checker_fence_regs_rd_cta_id[7><1] ,
         \warp_checker_fence_regs_rd_cta_id[7><0] ,
         \warp_checker_fence_regs_rd_cta_id[6><3] ,
         \warp_checker_fence_regs_rd_cta_id[6><2] ,
         \warp_checker_fence_regs_rd_cta_id[6><1] ,
         \warp_checker_fence_regs_rd_cta_id[6><0] ,
         \warp_checker_fence_regs_rd_cta_id[5><3] ,
         \warp_checker_fence_regs_rd_cta_id[5><2] ,
         \warp_checker_fence_regs_rd_cta_id[5><1] ,
         \warp_checker_fence_regs_rd_cta_id[5><0] ,
         \warp_checker_fence_regs_rd_cta_id[4><3] ,
         \warp_checker_fence_regs_rd_cta_id[4><2] ,
         \warp_checker_fence_regs_rd_cta_id[4><1] ,
         \warp_checker_fence_regs_rd_cta_id[4><0] ,
         \warp_checker_fence_regs_rd_cta_id[3><3] ,
         \warp_checker_fence_regs_rd_cta_id[3><2] ,
         \warp_checker_fence_regs_rd_cta_id[3><1] ,
         \warp_checker_fence_regs_rd_cta_id[3><0] ,
         \warp_checker_fence_regs_rd_cta_id[2><3] ,
         \warp_checker_fence_regs_rd_cta_id[2><2] ,
         \warp_checker_fence_regs_rd_cta_id[2><1] ,
         \warp_checker_fence_regs_rd_cta_id[2><0] ,
         \warp_checker_fence_regs_rd_cta_id[1><3] ,
         \warp_checker_fence_regs_rd_cta_id[1><2] ,
         \warp_checker_fence_regs_rd_cta_id[1><1] ,
         \warp_checker_fence_regs_rd_cta_id[1><0] ,
         \warp_checker_fence_regs_rd_cta_id[0><3] ,
         \warp_checker_fence_regs_rd_cta_id[0><2] ,
         \warp_checker_fence_regs_rd_cta_id[0><1] ,
         \warp_checker_fence_regs_rd_cta_id[0><0] ,
         \fence_regs_rd_cta_id[31><3] , \fence_regs_rd_cta_id[31><2] ,
         \fence_regs_rd_cta_id[31><1] , \fence_regs_rd_cta_id[31><0] ,
         \fence_regs_rd_cta_id[30><3] , \fence_regs_rd_cta_id[30><2] ,
         \fence_regs_rd_cta_id[30><1] , \fence_regs_rd_cta_id[30><0] ,
         \fence_regs_rd_cta_id[29><3] , \fence_regs_rd_cta_id[29><2] ,
         \fence_regs_rd_cta_id[29><1] , \fence_regs_rd_cta_id[29><0] ,
         \fence_regs_rd_cta_id[28><3] , \fence_regs_rd_cta_id[28><2] ,
         \fence_regs_rd_cta_id[28><1] , \fence_regs_rd_cta_id[28><0] ,
         \fence_regs_rd_cta_id[27><3] , \fence_regs_rd_cta_id[27><2] ,
         \fence_regs_rd_cta_id[27><1] , \fence_regs_rd_cta_id[27><0] ,
         \fence_regs_rd_cta_id[26><3] , \fence_regs_rd_cta_id[26><2] ,
         \fence_regs_rd_cta_id[26><1] , \fence_regs_rd_cta_id[26><0] ,
         \fence_regs_rd_cta_id[25><3] , \fence_regs_rd_cta_id[25><2] ,
         \fence_regs_rd_cta_id[25><1] , \fence_regs_rd_cta_id[25><0] ,
         \fence_regs_rd_cta_id[24><3] , \fence_regs_rd_cta_id[24><2] ,
         \fence_regs_rd_cta_id[24><1] , \fence_regs_rd_cta_id[24><0] ,
         \fence_regs_rd_cta_id[23><3] , \fence_regs_rd_cta_id[23><2] ,
         \fence_regs_rd_cta_id[23><1] , \fence_regs_rd_cta_id[23><0] ,
         \fence_regs_rd_cta_id[22><3] , \fence_regs_rd_cta_id[22><2] ,
         \fence_regs_rd_cta_id[22><1] , \fence_regs_rd_cta_id[22><0] ,
         \fence_regs_rd_cta_id[21><3] , \fence_regs_rd_cta_id[21><2] ,
         \fence_regs_rd_cta_id[21><1] , \fence_regs_rd_cta_id[21><0] ,
         \fence_regs_rd_cta_id[20><3] , \fence_regs_rd_cta_id[20><2] ,
         \fence_regs_rd_cta_id[20><1] , \fence_regs_rd_cta_id[20><0] ,
         \fence_regs_rd_cta_id[19><3] , \fence_regs_rd_cta_id[19><2] ,
         \fence_regs_rd_cta_id[19><1] , \fence_regs_rd_cta_id[19><0] ,
         \fence_regs_rd_cta_id[18><3] , \fence_regs_rd_cta_id[18><2] ,
         \fence_regs_rd_cta_id[18><1] , \fence_regs_rd_cta_id[18><0] ,
         \fence_regs_rd_cta_id[17><3] , \fence_regs_rd_cta_id[17><2] ,
         \fence_regs_rd_cta_id[17><1] , \fence_regs_rd_cta_id[17><0] ,
         \fence_regs_rd_cta_id[16><3] , \fence_regs_rd_cta_id[16><2] ,
         \fence_regs_rd_cta_id[16><1] , \fence_regs_rd_cta_id[16><0] ,
         \fence_regs_rd_cta_id[15><3] , \fence_regs_rd_cta_id[15><2] ,
         \fence_regs_rd_cta_id[15><1] , \fence_regs_rd_cta_id[15><0] ,
         \fence_regs_rd_cta_id[14><3] , \fence_regs_rd_cta_id[14><2] ,
         \fence_regs_rd_cta_id[14><1] , \fence_regs_rd_cta_id[14><0] ,
         \fence_regs_rd_cta_id[13><3] , \fence_regs_rd_cta_id[13><2] ,
         \fence_regs_rd_cta_id[13><1] , \fence_regs_rd_cta_id[13><0] ,
         \fence_regs_rd_cta_id[12><3] , \fence_regs_rd_cta_id[12><2] ,
         \fence_regs_rd_cta_id[12><1] , \fence_regs_rd_cta_id[12><0] ,
         \fence_regs_rd_cta_id[11><3] , \fence_regs_rd_cta_id[11><2] ,
         \fence_regs_rd_cta_id[11><1] , \fence_regs_rd_cta_id[11><0] ,
         \fence_regs_rd_cta_id[10><3] , \fence_regs_rd_cta_id[10><2] ,
         \fence_regs_rd_cta_id[10><1] , \fence_regs_rd_cta_id[10><0] ,
         \fence_regs_rd_cta_id[9><3] , \fence_regs_rd_cta_id[9><2] ,
         \fence_regs_rd_cta_id[9><1] , \fence_regs_rd_cta_id[9><0] ,
         \fence_regs_rd_cta_id[8><3] , \fence_regs_rd_cta_id[8><2] ,
         \fence_regs_rd_cta_id[8><1] , \fence_regs_rd_cta_id[8><0] ,
         \fence_regs_rd_cta_id[7><3] , \fence_regs_rd_cta_id[7><2] ,
         \fence_regs_rd_cta_id[7><1] , \fence_regs_rd_cta_id[7><0] ,
         \fence_regs_rd_cta_id[6><3] , \fence_regs_rd_cta_id[6><2] ,
         \fence_regs_rd_cta_id[6><1] , \fence_regs_rd_cta_id[6><0] ,
         \fence_regs_rd_cta_id[5><3] , \fence_regs_rd_cta_id[5><2] ,
         \fence_regs_rd_cta_id[5><1] , \fence_regs_rd_cta_id[5><0] ,
         \fence_regs_rd_cta_id[4><3] , \fence_regs_rd_cta_id[4><2] ,
         \fence_regs_rd_cta_id[4><1] , \fence_regs_rd_cta_id[4><0] ,
         \fence_regs_rd_cta_id[3><3] , \fence_regs_rd_cta_id[3><2] ,
         \fence_regs_rd_cta_id[3><1] , \fence_regs_rd_cta_id[3><0] ,
         \fence_regs_rd_cta_id[2><3] , \fence_regs_rd_cta_id[2><2] ,
         \fence_regs_rd_cta_id[2><1] , \fence_regs_rd_cta_id[2><0] ,
         \fence_regs_rd_cta_id[1><3] , \fence_regs_rd_cta_id[1><2] ,
         \fence_regs_rd_cta_id[1><1] , \fence_regs_rd_cta_id[1><0] ,
         \fence_regs_rd_cta_id[0><3] , \fence_regs_rd_cta_id[0><2] ,
         \fence_regs_rd_cta_id[0><1] , \fence_regs_rd_cta_id[0><0] ,
         \fence_regs_wr_cta_id[31><3] , \fence_regs_wr_cta_id[31><2] ,
         \fence_regs_wr_cta_id[31><1] , \fence_regs_wr_cta_id[31><0] ,
         \fence_regs_wr_cta_id[30><3] , \fence_regs_wr_cta_id[30><2] ,
         \fence_regs_wr_cta_id[30><1] , \fence_regs_wr_cta_id[30><0] ,
         \fence_regs_wr_cta_id[29><3] , \fence_regs_wr_cta_id[29><2] ,
         \fence_regs_wr_cta_id[29><1] , \fence_regs_wr_cta_id[29><0] ,
         \fence_regs_wr_cta_id[28><3] , \fence_regs_wr_cta_id[28><2] ,
         \fence_regs_wr_cta_id[28><1] , \fence_regs_wr_cta_id[28><0] ,
         \fence_regs_wr_cta_id[27><3] , \fence_regs_wr_cta_id[27><2] ,
         \fence_regs_wr_cta_id[27><1] , \fence_regs_wr_cta_id[27><0] ,
         \fence_regs_wr_cta_id[26><3] , \fence_regs_wr_cta_id[26><2] ,
         \fence_regs_wr_cta_id[26><1] , \fence_regs_wr_cta_id[26><0] ,
         \fence_regs_wr_cta_id[25><3] , \fence_regs_wr_cta_id[25><2] ,
         \fence_regs_wr_cta_id[25><1] , \fence_regs_wr_cta_id[25><0] ,
         \fence_regs_wr_cta_id[24><3] , \fence_regs_wr_cta_id[24><2] ,
         \fence_regs_wr_cta_id[24><1] , \fence_regs_wr_cta_id[24><0] ,
         \fence_regs_wr_cta_id[23><3] , \fence_regs_wr_cta_id[23><2] ,
         \fence_regs_wr_cta_id[23><1] , \fence_regs_wr_cta_id[23><0] ,
         \fence_regs_wr_cta_id[22><3] , \fence_regs_wr_cta_id[22><2] ,
         \fence_regs_wr_cta_id[22><1] , \fence_regs_wr_cta_id[22><0] ,
         \fence_regs_wr_cta_id[21><3] , \fence_regs_wr_cta_id[21><2] ,
         \fence_regs_wr_cta_id[21><1] , \fence_regs_wr_cta_id[21><0] ,
         \fence_regs_wr_cta_id[20><3] , \fence_regs_wr_cta_id[20><2] ,
         \fence_regs_wr_cta_id[20><1] , \fence_regs_wr_cta_id[20><0] ,
         \fence_regs_wr_cta_id[19><3] , \fence_regs_wr_cta_id[19><2] ,
         \fence_regs_wr_cta_id[19><1] , \fence_regs_wr_cta_id[19><0] ,
         \fence_regs_wr_cta_id[18><3] , \fence_regs_wr_cta_id[18><2] ,
         \fence_regs_wr_cta_id[18><1] , \fence_regs_wr_cta_id[18><0] ,
         \fence_regs_wr_cta_id[17><3] , \fence_regs_wr_cta_id[17><2] ,
         \fence_regs_wr_cta_id[17><1] , \fence_regs_wr_cta_id[17><0] ,
         \fence_regs_wr_cta_id[16><3] , \fence_regs_wr_cta_id[16><2] ,
         \fence_regs_wr_cta_id[16><1] , \fence_regs_wr_cta_id[16><0] ,
         \fence_regs_wr_cta_id[15><3] , \fence_regs_wr_cta_id[15><2] ,
         \fence_regs_wr_cta_id[15><1] , \fence_regs_wr_cta_id[15><0] ,
         \fence_regs_wr_cta_id[14><3] , \fence_regs_wr_cta_id[14><2] ,
         \fence_regs_wr_cta_id[14><1] , \fence_regs_wr_cta_id[14><0] ,
         \fence_regs_wr_cta_id[13><3] , \fence_regs_wr_cta_id[13><2] ,
         \fence_regs_wr_cta_id[13><1] , \fence_regs_wr_cta_id[13><0] ,
         \fence_regs_wr_cta_id[12><3] , \fence_regs_wr_cta_id[12><2] ,
         \fence_regs_wr_cta_id[12><1] , \fence_regs_wr_cta_id[12><0] ,
         \fence_regs_wr_cta_id[11><3] , \fence_regs_wr_cta_id[11><2] ,
         \fence_regs_wr_cta_id[11><1] , \fence_regs_wr_cta_id[11><0] ,
         \fence_regs_wr_cta_id[10><3] , \fence_regs_wr_cta_id[10><2] ,
         \fence_regs_wr_cta_id[10><1] , \fence_regs_wr_cta_id[10><0] ,
         \fence_regs_wr_cta_id[9><3] , \fence_regs_wr_cta_id[9><2] ,
         \fence_regs_wr_cta_id[9><1] , \fence_regs_wr_cta_id[9><0] ,
         \fence_regs_wr_cta_id[8><3] , \fence_regs_wr_cta_id[8><2] ,
         \fence_regs_wr_cta_id[8><1] , \fence_regs_wr_cta_id[8><0] ,
         \fence_regs_wr_cta_id[7><3] , \fence_regs_wr_cta_id[7><2] ,
         \fence_regs_wr_cta_id[7><1] , \fence_regs_wr_cta_id[7><0] ,
         \fence_regs_wr_cta_id[6><3] , \fence_regs_wr_cta_id[6><2] ,
         \fence_regs_wr_cta_id[6><1] , \fence_regs_wr_cta_id[6><0] ,
         \fence_regs_wr_cta_id[5><3] , \fence_regs_wr_cta_id[5><2] ,
         \fence_regs_wr_cta_id[5><1] , \fence_regs_wr_cta_id[5><0] ,
         \fence_regs_wr_cta_id[4><3] , \fence_regs_wr_cta_id[4><2] ,
         \fence_regs_wr_cta_id[4><1] , \fence_regs_wr_cta_id[4><0] ,
         \fence_regs_wr_cta_id[3><3] , \fence_regs_wr_cta_id[3><2] ,
         \fence_regs_wr_cta_id[3><1] , \fence_regs_wr_cta_id[3><0] ,
         \fence_regs_wr_cta_id[2><3] , \fence_regs_wr_cta_id[2><2] ,
         \fence_regs_wr_cta_id[2><1] , \fence_regs_wr_cta_id[2><0] ,
         \fence_regs_wr_cta_id[1><3] , \fence_regs_wr_cta_id[1><2] ,
         \fence_regs_wr_cta_id[1><1] , \fence_regs_wr_cta_id[1><0] ,
         \fence_regs_wr_cta_id[0><3] , \fence_regs_wr_cta_id[0><2] ,
         \fence_regs_wr_cta_id[0><1] , \fence_regs_wr_cta_id[0><0] , n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n208, n211, n212, n213, n214, n215, n345, n346, n347, n348, n349,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n209, n210, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261;
  wire   [4:0] warp_gen_pool_addr;
  wire   [127:0] warp_gen_pool_wr_data;
  wire   [4:0] warp_gen_state_addr;
  wire   [31:0] warp_gen_fence_regs_cta_id_ld;
  wire   [31:0] warp_gen_fence_regs_fence_en_ld;
  wire   [31:0] warps_done_mask_int;
  wire   [4:0] warp_sched_pool_addr;
  wire   [4:0] warp_sched_state_addr;
  wire   [4:0] warp_pool_addr_b;
  wire   [127:0] warp_pool_wr_data_b;
  wire   [4:0] warp_state_addr_b;
  wire   [1:0] warp_state_wr_data_b;
  wire   [31:0] warp_checker_fence_regs_wr_fence_en;
  wire   [31:0] warp_checker_fence_regs_fence_en_ld;
  wire   [31:0] warp_checker_fence_regs_rd_fence_en;
  wire   [127:0] warp_pool_rd_data_a;
  wire   [1:0] warp_state_rd_data_a;
  wire   [31:0] fence_regs_rd_fence_en;
  wire   [31:0] fence_regs_cta_id_ld;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42;

  warp_generator uWarpGenerator ( .clk_in(clk_in), 
        .host_reset(n248), .en(warp_generator_en), .num_blocks_in(
        num_blocks_in), .warps_per_block_in(warps_per_block_in), 
        .shmem_base_addr_in(shared_mem_base_addr_in), .shmem_size_in(
        shared_mem_size_in), .gprs_size_in(gprs_size_in), .warp_pool_addr_out(
        warp_gen_pool_addr), .warp_pool_wr_en_out(warp_gen_pool_wr_en), 
        .warp_pool_wr_data_out({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, warp_gen_pool_wr_data[123:97], 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, warp_gen_pool_wr_data[63:0]}), 
        .warp_state_addr_out(warp_gen_state_addr), .warp_state_wr_en_out(
        warp_gen_state_wr_en), .fence_regs_cta_id_out({
        \warp_gen_fence_regs_wr_cta_id[31><3] , 
        \warp_gen_fence_regs_wr_cta_id[31><2] , 
        \warp_gen_fence_regs_wr_cta_id[31><1] , 
        \warp_gen_fence_regs_wr_cta_id[31><0] , 
        \warp_gen_fence_regs_wr_cta_id[30><3] , 
        \warp_gen_fence_regs_wr_cta_id[30><2] , 
        \warp_gen_fence_regs_wr_cta_id[30><1] , 
        \warp_gen_fence_regs_wr_cta_id[30><0] , 
        \warp_gen_fence_regs_wr_cta_id[29><3] , 
        \warp_gen_fence_regs_wr_cta_id[29><2] , 
        \warp_gen_fence_regs_wr_cta_id[29><1] , 
        \warp_gen_fence_regs_wr_cta_id[29><0] , 
        \warp_gen_fence_regs_wr_cta_id[28><3] , 
        \warp_gen_fence_regs_wr_cta_id[28><2] , 
        \warp_gen_fence_regs_wr_cta_id[28><1] , 
        \warp_gen_fence_regs_wr_cta_id[28><0] , 
        \warp_gen_fence_regs_wr_cta_id[27><3] , 
        \warp_gen_fence_regs_wr_cta_id[27><2] , 
        \warp_gen_fence_regs_wr_cta_id[27><1] , 
        \warp_gen_fence_regs_wr_cta_id[27><0] , 
        \warp_gen_fence_regs_wr_cta_id[26><3] , 
        \warp_gen_fence_regs_wr_cta_id[26><2] , 
        \warp_gen_fence_regs_wr_cta_id[26><1] , 
        \warp_gen_fence_regs_wr_cta_id[26><0] , 
        \warp_gen_fence_regs_wr_cta_id[25><3] , 
        \warp_gen_fence_regs_wr_cta_id[25><2] , 
        \warp_gen_fence_regs_wr_cta_id[25><1] , 
        \warp_gen_fence_regs_wr_cta_id[25><0] , 
        \warp_gen_fence_regs_wr_cta_id[24><3] , 
        \warp_gen_fence_regs_wr_cta_id[24><2] , 
        \warp_gen_fence_regs_wr_cta_id[24><1] , 
        \warp_gen_fence_regs_wr_cta_id[24><0] , 
        \warp_gen_fence_regs_wr_cta_id[23><3] , 
        \warp_gen_fence_regs_wr_cta_id[23><2] , 
        \warp_gen_fence_regs_wr_cta_id[23><1] , 
        \warp_gen_fence_regs_wr_cta_id[23><0] , 
        \warp_gen_fence_regs_wr_cta_id[22><3] , 
        \warp_gen_fence_regs_wr_cta_id[22><2] , 
        \warp_gen_fence_regs_wr_cta_id[22><1] , 
        \warp_gen_fence_regs_wr_cta_id[22><0] , 
        \warp_gen_fence_regs_wr_cta_id[21><3] , 
        \warp_gen_fence_regs_wr_cta_id[21><2] , 
        \warp_gen_fence_regs_wr_cta_id[21><1] , 
        \warp_gen_fence_regs_wr_cta_id[21><0] , 
        \warp_gen_fence_regs_wr_cta_id[20><3] , 
        \warp_gen_fence_regs_wr_cta_id[20><2] , 
        \warp_gen_fence_regs_wr_cta_id[20><1] , 
        \warp_gen_fence_regs_wr_cta_id[20><0] , 
        \warp_gen_fence_regs_wr_cta_id[19><3] , 
        \warp_gen_fence_regs_wr_cta_id[19><2] , 
        \warp_gen_fence_regs_wr_cta_id[19><1] , 
        \warp_gen_fence_regs_wr_cta_id[19><0] , 
        \warp_gen_fence_regs_wr_cta_id[18><3] , 
        \warp_gen_fence_regs_wr_cta_id[18><2] , 
        \warp_gen_fence_regs_wr_cta_id[18><1] , 
        \warp_gen_fence_regs_wr_cta_id[18><0] , 
        \warp_gen_fence_regs_wr_cta_id[17><3] , 
        \warp_gen_fence_regs_wr_cta_id[17><2] , 
        \warp_gen_fence_regs_wr_cta_id[17><1] , 
        \warp_gen_fence_regs_wr_cta_id[17><0] , 
        \warp_gen_fence_regs_wr_cta_id[16><3] , 
        \warp_gen_fence_regs_wr_cta_id[16><2] , 
        \warp_gen_fence_regs_wr_cta_id[16><1] , 
        \warp_gen_fence_regs_wr_cta_id[16><0] , 
        \warp_gen_fence_regs_wr_cta_id[15><3] , 
        \warp_gen_fence_regs_wr_cta_id[15><2] , 
        \warp_gen_fence_regs_wr_cta_id[15><1] , 
        \warp_gen_fence_regs_wr_cta_id[15><0] , 
        \warp_gen_fence_regs_wr_cta_id[14><3] , 
        \warp_gen_fence_regs_wr_cta_id[14><2] , 
        \warp_gen_fence_regs_wr_cta_id[14><1] , 
        \warp_gen_fence_regs_wr_cta_id[14><0] , 
        \warp_gen_fence_regs_wr_cta_id[13><3] , 
        \warp_gen_fence_regs_wr_cta_id[13><2] , 
        \warp_gen_fence_regs_wr_cta_id[13><1] , 
        \warp_gen_fence_regs_wr_cta_id[13><0] , 
        \warp_gen_fence_regs_wr_cta_id[12><3] , 
        \warp_gen_fence_regs_wr_cta_id[12><2] , 
        \warp_gen_fence_regs_wr_cta_id[12><1] , 
        \warp_gen_fence_regs_wr_cta_id[12><0] , 
        \warp_gen_fence_regs_wr_cta_id[11><3] , 
        \warp_gen_fence_regs_wr_cta_id[11><2] , 
        \warp_gen_fence_regs_wr_cta_id[11><1] , 
        \warp_gen_fence_regs_wr_cta_id[11><0] , 
        \warp_gen_fence_regs_wr_cta_id[10><3] , 
        \warp_gen_fence_regs_wr_cta_id[10><2] , 
        \warp_gen_fence_regs_wr_cta_id[10><1] , 
        \warp_gen_fence_regs_wr_cta_id[10><0] , 
        \warp_gen_fence_regs_wr_cta_id[9><3] , 
        \warp_gen_fence_regs_wr_cta_id[9><2] , 
        \warp_gen_fence_regs_wr_cta_id[9><1] , 
        \warp_gen_fence_regs_wr_cta_id[9><0] , 
        \warp_gen_fence_regs_wr_cta_id[8><3] , 
        \warp_gen_fence_regs_wr_cta_id[8><2] , 
        \warp_gen_fence_regs_wr_cta_id[8><1] , 
        \warp_gen_fence_regs_wr_cta_id[8><0] , 
        \warp_gen_fence_regs_wr_cta_id[7><3] , 
        \warp_gen_fence_regs_wr_cta_id[7><2] , 
        \warp_gen_fence_regs_wr_cta_id[7><1] , 
        \warp_gen_fence_regs_wr_cta_id[7><0] , 
        \warp_gen_fence_regs_wr_cta_id[6><3] , 
        \warp_gen_fence_regs_wr_cta_id[6><2] , 
        \warp_gen_fence_regs_wr_cta_id[6><1] , 
        \warp_gen_fence_regs_wr_cta_id[6><0] , 
        \warp_gen_fence_regs_wr_cta_id[5><3] , 
        \warp_gen_fence_regs_wr_cta_id[5><2] , 
        \warp_gen_fence_regs_wr_cta_id[5><1] , 
        \warp_gen_fence_regs_wr_cta_id[5><0] , 
        \warp_gen_fence_regs_wr_cta_id[4><3] , 
        \warp_gen_fence_regs_wr_cta_id[4><2] , 
        \warp_gen_fence_regs_wr_cta_id[4><1] , 
        \warp_gen_fence_regs_wr_cta_id[4><0] , 
        \warp_gen_fence_regs_wr_cta_id[3><3] , 
        \warp_gen_fence_regs_wr_cta_id[3><2] , 
        \warp_gen_fence_regs_wr_cta_id[3><1] , 
        \warp_gen_fence_regs_wr_cta_id[3><0] , 
        \warp_gen_fence_regs_wr_cta_id[2><3] , 
        \warp_gen_fence_regs_wr_cta_id[2><2] , 
        \warp_gen_fence_regs_wr_cta_id[2><1] , 
        \warp_gen_fence_regs_wr_cta_id[2><0] , 
        \warp_gen_fence_regs_wr_cta_id[1><3] , 
        \warp_gen_fence_regs_wr_cta_id[1><2] , 
        \warp_gen_fence_regs_wr_cta_id[1><1] , 
        \warp_gen_fence_regs_wr_cta_id[1><0] , 
        \warp_gen_fence_regs_wr_cta_id[0><3] , 
        \warp_gen_fence_regs_wr_cta_id[0><2] , 
        \warp_gen_fence_regs_wr_cta_id[0><1] , 
        \warp_gen_fence_regs_wr_cta_id[0><0] }), .fence_regs_cta_id_ld(
        warp_gen_fence_regs_cta_id_ld), .fence_regs_fence_en_ld(
        warp_gen_fence_regs_fence_en_ld), .num_warps_out(num_warps_out), 
        .warp_gen_done(warp_generator_done) );
		
  warp_scheduler uWarpScheduler ( .clk_in(clk_in), 
        .host_reset(n248), .reset(n164), .pipeline_stall_in(pipeline_stall_in), 
        .num_blocks_in(num_blocks_in), .num_warps_in(num_warps_out), 
        .gprs_size_in(gprs_size_in), .warps_done_mask_in(warps_done_mask_int), 
        .warp_pool_addr_out(warp_sched_pool_addr), .warp_pool_rd_data_in(
        warp_pool_rd_data_a), .warp_state_addr_out(warp_sched_state_addr), 
        .warp_state_wr_en_out(warp_sched_state_wr_en), 
        .warp_state_wr_data_out({SYNOPSYS_UNCONNECTED__37, 
        \warp_sched_state_wr_data[0] }), .warp_state_rd_data_in(
        warp_state_rd_data_a), .program_cntr_out(program_cntr_out), 
        .warp_id_out(warp_id_out), .warp_lane_id_out(warp_lane_id_out), 
        .cta_id_out(cta_id_out), .initial_mask_out(initial_mask_out), 
        .current_mask_out(current_mask_out), .shmem_base_addr_out(
        shmem_base_addr_out), .gprs_size_out(gprs_size_out), 
        .gprs_base_addr_out(gprs_base_addr_out), .done(warp_scheduler_done), 
        .pipeline_warpunit_done(pipeline_warpunit_done), .fetch_en(fetch_en)
         );
  warp_checker uWarpChecker ( .clk_in(clk_in), .host_reset(
        n249), .reset(n164), .en(pipeline_write_done), .warp_id_in(warp_id_in), 
        .warp_lane_id_in(warp_lane_id_in), .cta_id_in(cta_id_in), 
        .initial_mask_in(initial_mask_in), .current_mask_in(current_mask_in), 
        .shmem_base_addr_in(shmem_base_addr_in), .gprs_base_addr_in(
        gprs_base_addr_in), .next_pc_in(next_pc_in), .warp_state_in(
        warp_state_in), .warps_per_block_in(warps_per_block_in), 
        .warp_pool_addr_out(warp_pool_addr_b), .warp_pool_wr_en_out(
        warp_pool_wr_en_b), .warp_pool_wr_data_out({SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, warp_pool_wr_data_b[123:97], 
        SYNOPSYS_UNCONNECTED__42, warp_pool_wr_data_b[95:0]}), 
        .warp_state_addr_out(warp_state_addr_b), .warp_state_wr_en_out(
        warp_state_wr_en_b), .warp_state_wr_data_out(warp_state_wr_data_b), 
        .fence_regs_fence_en_out(warp_checker_fence_regs_wr_fence_en), 
        .fence_regs_fence_en_ld(warp_checker_fence_regs_fence_en_ld), 
        .fence_regs_cta_id_in({\warp_checker_fence_regs_rd_cta_id[31><3] , 
        \warp_checker_fence_regs_rd_cta_id[31><2] , 
        \warp_checker_fence_regs_rd_cta_id[31><1] , 
        \warp_checker_fence_regs_rd_cta_id[31><0] , 
        \warp_checker_fence_regs_rd_cta_id[30><3] , 
        \warp_checker_fence_regs_rd_cta_id[30><2] , 
        \warp_checker_fence_regs_rd_cta_id[30><1] , 
        \warp_checker_fence_regs_rd_cta_id[30><0] , 
        \warp_checker_fence_regs_rd_cta_id[29><3] , 
        \warp_checker_fence_regs_rd_cta_id[29><2] , 
        \warp_checker_fence_regs_rd_cta_id[29><1] , 
        \warp_checker_fence_regs_rd_cta_id[29><0] , 
        \warp_checker_fence_regs_rd_cta_id[28><3] , 
        \warp_checker_fence_regs_rd_cta_id[28><2] , 
        \warp_checker_fence_regs_rd_cta_id[28><1] , 
        \warp_checker_fence_regs_rd_cta_id[28><0] , 
        \warp_checker_fence_regs_rd_cta_id[27><3] , 
        \warp_checker_fence_regs_rd_cta_id[27><2] , 
        \warp_checker_fence_regs_rd_cta_id[27><1] , 
        \warp_checker_fence_regs_rd_cta_id[27><0] , 
        \warp_checker_fence_regs_rd_cta_id[26><3] , 
        \warp_checker_fence_regs_rd_cta_id[26><2] , 
        \warp_checker_fence_regs_rd_cta_id[26><1] , 
        \warp_checker_fence_regs_rd_cta_id[26><0] , 
        \warp_checker_fence_regs_rd_cta_id[25><3] , 
        \warp_checker_fence_regs_rd_cta_id[25><2] , 
        \warp_checker_fence_regs_rd_cta_id[25><1] , 
        \warp_checker_fence_regs_rd_cta_id[25><0] , 
        \warp_checker_fence_regs_rd_cta_id[24><3] , 
        \warp_checker_fence_regs_rd_cta_id[24><2] , 
        \warp_checker_fence_regs_rd_cta_id[24><1] , 
        \warp_checker_fence_regs_rd_cta_id[24><0] , 
        \warp_checker_fence_regs_rd_cta_id[23><3] , 
        \warp_checker_fence_regs_rd_cta_id[23><2] , 
        \warp_checker_fence_regs_rd_cta_id[23><1] , 
        \warp_checker_fence_regs_rd_cta_id[23><0] , 
        \warp_checker_fence_regs_rd_cta_id[22><3] , 
        \warp_checker_fence_regs_rd_cta_id[22><2] , 
        \warp_checker_fence_regs_rd_cta_id[22><1] , 
        \warp_checker_fence_regs_rd_cta_id[22><0] , 
        \warp_checker_fence_regs_rd_cta_id[21><3] , 
        \warp_checker_fence_regs_rd_cta_id[21><2] , 
        \warp_checker_fence_regs_rd_cta_id[21><1] , 
        \warp_checker_fence_regs_rd_cta_id[21><0] , 
        \warp_checker_fence_regs_rd_cta_id[20><3] , 
        \warp_checker_fence_regs_rd_cta_id[20><2] , 
        \warp_checker_fence_regs_rd_cta_id[20><1] , 
        \warp_checker_fence_regs_rd_cta_id[20><0] , 
        \warp_checker_fence_regs_rd_cta_id[19><3] , 
        \warp_checker_fence_regs_rd_cta_id[19><2] , 
        \warp_checker_fence_regs_rd_cta_id[19><1] , 
        \warp_checker_fence_regs_rd_cta_id[19><0] , 
        \warp_checker_fence_regs_rd_cta_id[18><3] , 
        \warp_checker_fence_regs_rd_cta_id[18><2] , 
        \warp_checker_fence_regs_rd_cta_id[18><1] , 
        \warp_checker_fence_regs_rd_cta_id[18><0] , 
        \warp_checker_fence_regs_rd_cta_id[17><3] , 
        \warp_checker_fence_regs_rd_cta_id[17><2] , 
        \warp_checker_fence_regs_rd_cta_id[17><1] , 
        \warp_checker_fence_regs_rd_cta_id[17><0] , 
        \warp_checker_fence_regs_rd_cta_id[16><3] , 
        \warp_checker_fence_regs_rd_cta_id[16><2] , 
        \warp_checker_fence_regs_rd_cta_id[16><1] , 
        \warp_checker_fence_regs_rd_cta_id[16><0] , 
        \warp_checker_fence_regs_rd_cta_id[15><3] , 
        \warp_checker_fence_regs_rd_cta_id[15><2] , 
        \warp_checker_fence_regs_rd_cta_id[15><1] , 
        \warp_checker_fence_regs_rd_cta_id[15><0] , 
        \warp_checker_fence_regs_rd_cta_id[14><3] , 
        \warp_checker_fence_regs_rd_cta_id[14><2] , 
        \warp_checker_fence_regs_rd_cta_id[14><1] , 
        \warp_checker_fence_regs_rd_cta_id[14><0] , 
        \warp_checker_fence_regs_rd_cta_id[13><3] , 
        \warp_checker_fence_regs_rd_cta_id[13><2] , 
        \warp_checker_fence_regs_rd_cta_id[13><1] , 
        \warp_checker_fence_regs_rd_cta_id[13><0] , 
        \warp_checker_fence_regs_rd_cta_id[12><3] , 
        \warp_checker_fence_regs_rd_cta_id[12><2] , 
        \warp_checker_fence_regs_rd_cta_id[12><1] , 
        \warp_checker_fence_regs_rd_cta_id[12><0] , 
        \warp_checker_fence_regs_rd_cta_id[11><3] , 
        \warp_checker_fence_regs_rd_cta_id[11><2] , 
        \warp_checker_fence_regs_rd_cta_id[11><1] , 
        \warp_checker_fence_regs_rd_cta_id[11><0] , 
        \warp_checker_fence_regs_rd_cta_id[10><3] , 
        \warp_checker_fence_regs_rd_cta_id[10><2] , 
        \warp_checker_fence_regs_rd_cta_id[10><1] , 
        \warp_checker_fence_regs_rd_cta_id[10><0] , 
        \warp_checker_fence_regs_rd_cta_id[9><3] , 
        \warp_checker_fence_regs_rd_cta_id[9><2] , 
        \warp_checker_fence_regs_rd_cta_id[9><1] , 
        \warp_checker_fence_regs_rd_cta_id[9><0] , 
        \warp_checker_fence_regs_rd_cta_id[8><3] , 
        \warp_checker_fence_regs_rd_cta_id[8><2] , 
        \warp_checker_fence_regs_rd_cta_id[8><1] , 
        \warp_checker_fence_regs_rd_cta_id[8><0] , 
        \warp_checker_fence_regs_rd_cta_id[7><3] , 
        \warp_checker_fence_regs_rd_cta_id[7><2] , 
        \warp_checker_fence_regs_rd_cta_id[7><1] , 
        \warp_checker_fence_regs_rd_cta_id[7><0] , 
        \warp_checker_fence_regs_rd_cta_id[6><3] , 
        \warp_checker_fence_regs_rd_cta_id[6><2] , 
        \warp_checker_fence_regs_rd_cta_id[6><1] , 
        \warp_checker_fence_regs_rd_cta_id[6><0] , 
        \warp_checker_fence_regs_rd_cta_id[5><3] , 
        \warp_checker_fence_regs_rd_cta_id[5><2] , 
        \warp_checker_fence_regs_rd_cta_id[5><1] , 
        \warp_checker_fence_regs_rd_cta_id[5><0] , 
        \warp_checker_fence_regs_rd_cta_id[4><3] , 
        \warp_checker_fence_regs_rd_cta_id[4><2] , 
        \warp_checker_fence_regs_rd_cta_id[4><1] , 
        \warp_checker_fence_regs_rd_cta_id[4><0] , 
        \warp_checker_fence_regs_rd_cta_id[3><3] , 
        \warp_checker_fence_regs_rd_cta_id[3><2] , 
        \warp_checker_fence_regs_rd_cta_id[3><1] , 
        \warp_checker_fence_regs_rd_cta_id[3><0] , 
        \warp_checker_fence_regs_rd_cta_id[2><3] , 
        \warp_checker_fence_regs_rd_cta_id[2><2] , 
        \warp_checker_fence_regs_rd_cta_id[2><1] , 
        \warp_checker_fence_regs_rd_cta_id[2><0] , 
        \warp_checker_fence_regs_rd_cta_id[1><3] , 
        \warp_checker_fence_regs_rd_cta_id[1><2] , 
        \warp_checker_fence_regs_rd_cta_id[1><1] , 
        \warp_checker_fence_regs_rd_cta_id[1><0] , 
        \warp_checker_fence_regs_rd_cta_id[0><3] , 
        \warp_checker_fence_regs_rd_cta_id[0><2] , 
        \warp_checker_fence_regs_rd_cta_id[0><1] , 
        \warp_checker_fence_regs_rd_cta_id[0><0] }), .fence_regs_fence_en_in(
        warp_checker_fence_regs_rd_fence_en), .warps_done_mask_out(
        warps_done_mask_int), .pipeline_stall_out(pipeline_stall_out) );
  dp_regfile_RAM_SIZE32_RAM_A_WIDTH5_RAM_D_WIDTH128_1 uWarpPoolMemory ( .clk(
        clk_in), .rst(n249), .addr_a({n259, n253, n255, n261, n257}), .din_a({
        1'b0, 1'b0, 1'b0, 1'b0, n88, n87, n86, n85, n84, n83, n82, n80, n79, 
        n78, n77, n76, n75, n74, n73, n72, n71, n70, n69, n68, n67, n66, n65, 
        n152, n151, n150, n149, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, n148, n147, n146, n145, n144, n143, n142, n141, n140, n139, n138, 
        n137, n104, n103, n102, n101, n100, n99, n98, n97, n96, n95, n94, n93, 
        n92, n91, n90, n136, n135, n134, n133, n132, n131, n130, n129, n128, 
        n127, n126, n125, n124, n123, n122, n121, n120, n119, n118, n117, n116, 
        n115, n114, n113, n112, n111, n110, n109, n108, n107, n106, n105, n156, 
        n155, n154, n153, n81}), .we_a(n89), .addr_b(warp_pool_addr_b), 
        .din_b({1'b0, 1'b0, 1'b0, 1'b0, warp_pool_wr_data_b[123:97], 1'b0, 
        warp_pool_wr_data_b[95:0]}), .we_b(warp_pool_wr_en_b), .dout_a(
        warp_pool_rd_data_a) );
  dp_regfile_RAM_SIZE32_RAM_A_WIDTH5_RAM_D_WIDTH2_1 uWarpStateMemory ( .clk(
        clk_in), .rst(n249), .addr_a({n258, n252, n254, n260, n256}), .din_a({
        1'b0, n157}), .we_a(n251), .addr_b(warp_state_addr_b), .din_b(
        warp_state_wr_data_b), .we_b(warp_state_wr_en_b), .dout_a(
        warp_state_rd_data_a) );
  fence_registers_1_0 uFenceRegisters_0 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[0><3] , \fence_regs_wr_cta_id[0><2] , 
        \fence_regs_wr_cta_id[0><1] , \fence_regs_wr_cta_id[0><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[0]), .fence_en_in(n55), .fence_en_ld(
        n1), .cta_id_out({\fence_regs_rd_cta_id[0><3] , 
        \fence_regs_rd_cta_id[0><2] , \fence_regs_rd_cta_id[0><1] , 
        \fence_regs_rd_cta_id[0><0] }), .fence_en_out(
        fence_regs_rd_fence_en[0]) );
  fence_registers_1_31 uFenceRegisters_1 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[1><3] , \fence_regs_wr_cta_id[1><2] , 
        \fence_regs_wr_cta_id[1><1] , \fence_regs_wr_cta_id[1><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[1]), .fence_en_in(n33), .fence_en_ld(
        n2), .cta_id_out({\fence_regs_rd_cta_id[1><3] , 
        \fence_regs_rd_cta_id[1><2] , \fence_regs_rd_cta_id[1><1] , 
        \fence_regs_rd_cta_id[1><0] }), .fence_en_out(
        fence_regs_rd_fence_en[1]) );
  fence_registers_1_30 uFenceRegisters_2 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[2><3] , \fence_regs_wr_cta_id[2><2] , 
        \fence_regs_wr_cta_id[2><1] , \fence_regs_wr_cta_id[2><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[2]), .fence_en_in(n34), .fence_en_ld(
        n3), .cta_id_out({\fence_regs_rd_cta_id[2><3] , 
        \fence_regs_rd_cta_id[2><2] , \fence_regs_rd_cta_id[2><1] , 
        \fence_regs_rd_cta_id[2><0] }), .fence_en_out(
        fence_regs_rd_fence_en[2]) );
  fence_registers_1_29 uFenceRegisters_3 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[3><3] , \fence_regs_wr_cta_id[3><2] , 
        \fence_regs_wr_cta_id[3><1] , \fence_regs_wr_cta_id[3><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[3]), .fence_en_in(n56), .fence_en_ld(
        n4), .cta_id_out({\fence_regs_rd_cta_id[3><3] , 
        \fence_regs_rd_cta_id[3><2] , \fence_regs_rd_cta_id[3><1] , 
        \fence_regs_rd_cta_id[3><0] }), .fence_en_out(
        fence_regs_rd_fence_en[3]) );
  fence_registers_1_28 uFenceRegisters_4 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[4><3] , \fence_regs_wr_cta_id[4><2] , 
        \fence_regs_wr_cta_id[4><1] , \fence_regs_wr_cta_id[4><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[4]), .fence_en_in(n35), .fence_en_ld(
        n5), .cta_id_out({\fence_regs_rd_cta_id[4><3] , 
        \fence_regs_rd_cta_id[4><2] , \fence_regs_rd_cta_id[4><1] , 
        \fence_regs_rd_cta_id[4><0] }), .fence_en_out(
        fence_regs_rd_fence_en[4]) );
  fence_registers_1_27 uFenceRegisters_5 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[5><3] , \fence_regs_wr_cta_id[5><2] , 
        \fence_regs_wr_cta_id[5><1] , \fence_regs_wr_cta_id[5><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[5]), .fence_en_in(n36), .fence_en_ld(
        n6), .cta_id_out({\fence_regs_rd_cta_id[5><3] , 
        \fence_regs_rd_cta_id[5><2] , \fence_regs_rd_cta_id[5><1] , 
        \fence_regs_rd_cta_id[5><0] }), .fence_en_out(
        fence_regs_rd_fence_en[5]) );
  fence_registers_1_26 uFenceRegisters_6 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[6><3] , \fence_regs_wr_cta_id[6><2] , 
        \fence_regs_wr_cta_id[6><1] , \fence_regs_wr_cta_id[6><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[6]), .fence_en_in(n37), .fence_en_ld(
        n7), .cta_id_out({\fence_regs_rd_cta_id[6><3] , 
        \fence_regs_rd_cta_id[6><2] , \fence_regs_rd_cta_id[6><1] , 
        \fence_regs_rd_cta_id[6><0] }), .fence_en_out(
        fence_regs_rd_fence_en[6]) );
  fence_registers_1_25 uFenceRegisters_7 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[7><3] , \fence_regs_wr_cta_id[7><2] , 
        \fence_regs_wr_cta_id[7><1] , \fence_regs_wr_cta_id[7><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[7]), .fence_en_in(n38), .fence_en_ld(
        n8), .cta_id_out({\fence_regs_rd_cta_id[7><3] , 
        \fence_regs_rd_cta_id[7><2] , \fence_regs_rd_cta_id[7><1] , 
        \fence_regs_rd_cta_id[7><0] }), .fence_en_out(
        fence_regs_rd_fence_en[7]) );
  fence_registers_1_24 uFenceRegisters_8 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[8><3] , \fence_regs_wr_cta_id[8><2] , 
        \fence_regs_wr_cta_id[8><1] , \fence_regs_wr_cta_id[8><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[8]), .fence_en_in(n39), .fence_en_ld(
        n9), .cta_id_out({\fence_regs_rd_cta_id[8><3] , 
        \fence_regs_rd_cta_id[8><2] , \fence_regs_rd_cta_id[8><1] , 
        \fence_regs_rd_cta_id[8><0] }), .fence_en_out(
        fence_regs_rd_fence_en[8]) );
  fence_registers_1_23 uFenceRegisters_9 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[9><3] , \fence_regs_wr_cta_id[9><2] , 
        \fence_regs_wr_cta_id[9><1] , \fence_regs_wr_cta_id[9><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[9]), .fence_en_in(n57), .fence_en_ld(
        n10), .cta_id_out({\fence_regs_rd_cta_id[9><3] , 
        \fence_regs_rd_cta_id[9><2] , \fence_regs_rd_cta_id[9><1] , 
        \fence_regs_rd_cta_id[9><0] }), .fence_en_out(
        fence_regs_rd_fence_en[9]) );
  fence_registers_1_22 uFenceRegisters_10 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[10><3] , 
        \fence_regs_wr_cta_id[10><2] , \fence_regs_wr_cta_id[10><1] , 
        \fence_regs_wr_cta_id[10><0] }), .cta_id_ld(fence_regs_cta_id_ld[10]), 
        .fence_en_in(n40), .fence_en_ld(n11), .cta_id_out({
        \fence_regs_rd_cta_id[10><3] , \fence_regs_rd_cta_id[10><2] , 
        \fence_regs_rd_cta_id[10><1] , \fence_regs_rd_cta_id[10><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[10]) );
  fence_registers_1_21 uFenceRegisters_11 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[11><3] , 
        \fence_regs_wr_cta_id[11><2] , \fence_regs_wr_cta_id[11><1] , 
        \fence_regs_wr_cta_id[11><0] }), .cta_id_ld(fence_regs_cta_id_ld[11]), 
        .fence_en_in(n41), .fence_en_ld(n12), .cta_id_out({
        \fence_regs_rd_cta_id[11><3] , \fence_regs_rd_cta_id[11><2] , 
        \fence_regs_rd_cta_id[11><1] , \fence_regs_rd_cta_id[11><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[11]) );
  fence_registers_1_20 uFenceRegisters_12 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[12><3] , 
        \fence_regs_wr_cta_id[12><2] , \fence_regs_wr_cta_id[12><1] , 
        \fence_regs_wr_cta_id[12><0] }), .cta_id_ld(fence_regs_cta_id_ld[12]), 
        .fence_en_in(n62), .fence_en_ld(n13), .cta_id_out({
        \fence_regs_rd_cta_id[12><3] , \fence_regs_rd_cta_id[12><2] , 
        \fence_regs_rd_cta_id[12><1] , \fence_regs_rd_cta_id[12><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[12]) );
  fence_registers_1_19 uFenceRegisters_13 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[13><3] , 
        \fence_regs_wr_cta_id[13><2] , \fence_regs_wr_cta_id[13><1] , 
        \fence_regs_wr_cta_id[13><0] }), .cta_id_ld(fence_regs_cta_id_ld[13]), 
        .fence_en_in(n42), .fence_en_ld(n14), .cta_id_out({
        \fence_regs_rd_cta_id[13><3] , \fence_regs_rd_cta_id[13><2] , 
        \fence_regs_rd_cta_id[13><1] , \fence_regs_rd_cta_id[13><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[13]) );
  fence_registers_1_18 uFenceRegisters_14 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[14><3] , 
        \fence_regs_wr_cta_id[14><2] , \fence_regs_wr_cta_id[14><1] , 
        \fence_regs_wr_cta_id[14><0] }), .cta_id_ld(fence_regs_cta_id_ld[14]), 
        .fence_en_in(n43), .fence_en_ld(n15), .cta_id_out({
        \fence_regs_rd_cta_id[14><3] , \fence_regs_rd_cta_id[14><2] , 
        \fence_regs_rd_cta_id[14><1] , \fence_regs_rd_cta_id[14><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[14]) );
  fence_registers_1_17 uFenceRegisters_15 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[15><3] , 
        \fence_regs_wr_cta_id[15><2] , \fence_regs_wr_cta_id[15><1] , 
        \fence_regs_wr_cta_id[15><0] }), .cta_id_ld(fence_regs_cta_id_ld[15]), 
        .fence_en_in(n58), .fence_en_ld(n16), .cta_id_out({
        \fence_regs_rd_cta_id[15><3] , \fence_regs_rd_cta_id[15><2] , 
        \fence_regs_rd_cta_id[15><1] , \fence_regs_rd_cta_id[15><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[15]) );
  fence_registers_1_16 uFenceRegisters_16 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[16><3] , 
        \fence_regs_wr_cta_id[16><2] , \fence_regs_wr_cta_id[16><1] , 
        \fence_regs_wr_cta_id[16><0] }), .cta_id_ld(fence_regs_cta_id_ld[16]), 
        .fence_en_in(n44), .fence_en_ld(n17), .cta_id_out({
        \fence_regs_rd_cta_id[16><3] , \fence_regs_rd_cta_id[16><2] , 
        \fence_regs_rd_cta_id[16><1] , \fence_regs_rd_cta_id[16><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[16]) );
  fence_registers_1_15 uFenceRegisters_17 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[17><3] , 
        \fence_regs_wr_cta_id[17><2] , \fence_regs_wr_cta_id[17><1] , 
        \fence_regs_wr_cta_id[17><0] }), .cta_id_ld(fence_regs_cta_id_ld[17]), 
        .fence_en_in(n63), .fence_en_ld(n18), .cta_id_out({
        \fence_regs_rd_cta_id[17><3] , \fence_regs_rd_cta_id[17><2] , 
        \fence_regs_rd_cta_id[17><1] , \fence_regs_rd_cta_id[17><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[17]) );
  fence_registers_1_14 uFenceRegisters_18 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[18><3] , 
        \fence_regs_wr_cta_id[18><2] , \fence_regs_wr_cta_id[18><1] , 
        \fence_regs_wr_cta_id[18><0] }), .cta_id_ld(fence_regs_cta_id_ld[18]), 
        .fence_en_in(n45), .fence_en_ld(n19), .cta_id_out({
        \fence_regs_rd_cta_id[18><3] , \fence_regs_rd_cta_id[18><2] , 
        \fence_regs_rd_cta_id[18><1] , \fence_regs_rd_cta_id[18><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[18]) );
  fence_registers_1_13 uFenceRegisters_19 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[19><3] , 
        \fence_regs_wr_cta_id[19><2] , \fence_regs_wr_cta_id[19><1] , 
        \fence_regs_wr_cta_id[19><0] }), .cta_id_ld(fence_regs_cta_id_ld[19]), 
        .fence_en_in(n46), .fence_en_ld(n20), .cta_id_out({
        \fence_regs_rd_cta_id[19><3] , \fence_regs_rd_cta_id[19><2] , 
        \fence_regs_rd_cta_id[19><1] , \fence_regs_rd_cta_id[19><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[19]) );
  fence_registers_1_12 uFenceRegisters_20 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[20><3] , 
        \fence_regs_wr_cta_id[20><2] , \fence_regs_wr_cta_id[20><1] , 
        \fence_regs_wr_cta_id[20><0] }), .cta_id_ld(fence_regs_cta_id_ld[20]), 
        .fence_en_in(n47), .fence_en_ld(n21), .cta_id_out({
        \fence_regs_rd_cta_id[20><3] , \fence_regs_rd_cta_id[20><2] , 
        \fence_regs_rd_cta_id[20><1] , \fence_regs_rd_cta_id[20><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[20]) );
  fence_registers_1_11 uFenceRegisters_21 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[21><3] , 
        \fence_regs_wr_cta_id[21><2] , \fence_regs_wr_cta_id[21><1] , 
        \fence_regs_wr_cta_id[21><0] }), .cta_id_ld(fence_regs_cta_id_ld[21]), 
        .fence_en_in(n48), .fence_en_ld(n22), .cta_id_out({
        \fence_regs_rd_cta_id[21><3] , \fence_regs_rd_cta_id[21><2] , 
        \fence_regs_rd_cta_id[21><1] , \fence_regs_rd_cta_id[21><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[21]) );
  fence_registers_1_10 uFenceRegisters_22 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[22><3] , 
        \fence_regs_wr_cta_id[22><2] , \fence_regs_wr_cta_id[22><1] , 
        \fence_regs_wr_cta_id[22><0] }), .cta_id_ld(fence_regs_cta_id_ld[22]), 
        .fence_en_in(n49), .fence_en_ld(n23), .cta_id_out({
        \fence_regs_rd_cta_id[22><3] , \fence_regs_rd_cta_id[22><2] , 
        \fence_regs_rd_cta_id[22><1] , \fence_regs_rd_cta_id[22><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[22]) );
  fence_registers_1_9 uFenceRegisters_23 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[23><3] , 
        \fence_regs_wr_cta_id[23><2] , \fence_regs_wr_cta_id[23><1] , 
        \fence_regs_wr_cta_id[23><0] }), .cta_id_ld(fence_regs_cta_id_ld[23]), 
        .fence_en_in(n50), .fence_en_ld(n24), .cta_id_out({
        \fence_regs_rd_cta_id[23><3] , \fence_regs_rd_cta_id[23><2] , 
        \fence_regs_rd_cta_id[23><1] , \fence_regs_rd_cta_id[23><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[23]) );
  fence_registers_1_8 uFenceRegisters_24 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[24><3] , 
        \fence_regs_wr_cta_id[24><2] , \fence_regs_wr_cta_id[24><1] , 
        \fence_regs_wr_cta_id[24><0] }), .cta_id_ld(fence_regs_cta_id_ld[24]), 
        .fence_en_in(n51), .fence_en_ld(n25), .cta_id_out({
        \fence_regs_rd_cta_id[24><3] , \fence_regs_rd_cta_id[24><2] , 
        \fence_regs_rd_cta_id[24><1] , \fence_regs_rd_cta_id[24><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[24]) );
  fence_registers_1_7 uFenceRegisters_25 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[25><3] , 
        \fence_regs_wr_cta_id[25><2] , \fence_regs_wr_cta_id[25><1] , 
        \fence_regs_wr_cta_id[25><0] }), .cta_id_ld(fence_regs_cta_id_ld[25]), 
        .fence_en_in(n52), .fence_en_ld(n26), .cta_id_out({
        \fence_regs_rd_cta_id[25><3] , \fence_regs_rd_cta_id[25><2] , 
        \fence_regs_rd_cta_id[25><1] , \fence_regs_rd_cta_id[25><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[25]) );
  fence_registers_1_6 uFenceRegisters_26 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[26><3] , 
        \fence_regs_wr_cta_id[26><2] , \fence_regs_wr_cta_id[26><1] , 
        \fence_regs_wr_cta_id[26><0] }), .cta_id_ld(fence_regs_cta_id_ld[26]), 
        .fence_en_in(n53), .fence_en_ld(n27), .cta_id_out({
        \fence_regs_rd_cta_id[26><3] , \fence_regs_rd_cta_id[26><2] , 
        \fence_regs_rd_cta_id[26><1] , \fence_regs_rd_cta_id[26><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[26]) );
  fence_registers_1_5 uFenceRegisters_27 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[27><3] , 
        \fence_regs_wr_cta_id[27><2] , \fence_regs_wr_cta_id[27><1] , 
        \fence_regs_wr_cta_id[27><0] }), .cta_id_ld(fence_regs_cta_id_ld[27]), 
        .fence_en_in(n54), .fence_en_ld(n28), .cta_id_out({
        \fence_regs_rd_cta_id[27><3] , \fence_regs_rd_cta_id[27><2] , 
        \fence_regs_rd_cta_id[27><1] , \fence_regs_rd_cta_id[27><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[27]) );
  fence_registers_1_4 uFenceRegisters_28 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[28><3] , 
        \fence_regs_wr_cta_id[28><2] , \fence_regs_wr_cta_id[28><1] , 
        \fence_regs_wr_cta_id[28><0] }), .cta_id_ld(fence_regs_cta_id_ld[28]), 
        .fence_en_in(n59), .fence_en_ld(n29), .cta_id_out({
        \fence_regs_rd_cta_id[28><3] , \fence_regs_rd_cta_id[28><2] , 
        \fence_regs_rd_cta_id[28><1] , \fence_regs_rd_cta_id[28><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[28]) );
  fence_registers_1_3 uFenceRegisters_29 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[29><3] , 
        \fence_regs_wr_cta_id[29><2] , \fence_regs_wr_cta_id[29><1] , 
        \fence_regs_wr_cta_id[29><0] }), .cta_id_ld(fence_regs_cta_id_ld[29]), 
        .fence_en_in(n60), .fence_en_ld(n30), .cta_id_out({
        \fence_regs_rd_cta_id[29><3] , \fence_regs_rd_cta_id[29><2] , 
        \fence_regs_rd_cta_id[29><1] , \fence_regs_rd_cta_id[29><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[29]) );
  fence_registers_1_2 uFenceRegisters_30 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[30><3] , 
        \fence_regs_wr_cta_id[30><2] , \fence_regs_wr_cta_id[30><1] , 
        \fence_regs_wr_cta_id[30><0] }), .cta_id_ld(fence_regs_cta_id_ld[30]), 
        .fence_en_in(n64), .fence_en_ld(n31), .cta_id_out({
        \fence_regs_rd_cta_id[30><3] , \fence_regs_rd_cta_id[30><2] , 
        \fence_regs_rd_cta_id[30><1] , \fence_regs_rd_cta_id[30><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[30]) );
  fence_registers_1_1 uFenceRegisters_31 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[31><3] , 
        \fence_regs_wr_cta_id[31><2] , \fence_regs_wr_cta_id[31><1] , 
        \fence_regs_wr_cta_id[31><0] }), .cta_id_ld(fence_regs_cta_id_ld[31]), 
        .fence_en_in(n61), .fence_en_ld(n32), .cta_id_out({
        \fence_regs_rd_cta_id[31><3] , \fence_regs_rd_cta_id[31><2] , 
        \fence_regs_rd_cta_id[31><1] , \fence_regs_rd_cta_id[31><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[31]) );
  AND2_X1 U3 ( .A1(warp_checker_fence_regs_wr_fence_en[1]), .A2(n221), .ZN(n33) );
  AND2_X1 U4 ( .A1(warp_checker_fence_regs_wr_fence_en[2]), .A2(n221), .ZN(n34) );
  AND2_X1 U5 ( .A1(warp_checker_fence_regs_wr_fence_en[4]), .A2(n222), .ZN(n35) );
  AND2_X1 U6 ( .A1(warp_checker_fence_regs_wr_fence_en[5]), .A2(n223), .ZN(n36) );
  AND2_X1 U7 ( .A1(warp_checker_fence_regs_wr_fence_en[6]), .A2(n223), .ZN(n37) );
  AND2_X1 U8 ( .A1(warp_checker_fence_regs_wr_fence_en[7]), .A2(n222), .ZN(n38) );
  AND2_X1 U9 ( .A1(warp_checker_fence_regs_wr_fence_en[8]), .A2(n222), .ZN(n39) );
  AND2_X1 U10 ( .A1(warp_checker_fence_regs_wr_fence_en[10]), .A2(n222), .ZN(
        n40) );
  AND2_X1 U11 ( .A1(warp_checker_fence_regs_wr_fence_en[11]), .A2(n222), .ZN(
        n41) );
  AND2_X1 U12 ( .A1(warp_checker_fence_regs_wr_fence_en[13]), .A2(n222), .ZN(
        n42) );
  AND2_X1 U13 ( .A1(warp_checker_fence_regs_wr_fence_en[14]), .A2(n222), .ZN(
        n43) );
  AND2_X1 U14 ( .A1(warp_checker_fence_regs_wr_fence_en[16]), .A2(n223), .ZN(
        n44) );
  AND2_X1 U15 ( .A1(warp_checker_fence_regs_wr_fence_en[18]), .A2(n225), .ZN(
        n45) );
  AND2_X1 U16 ( .A1(warp_checker_fence_regs_wr_fence_en[19]), .A2(n225), .ZN(
        n46) );
  AND2_X1 U17 ( .A1(warp_checker_fence_regs_wr_fence_en[20]), .A2(n223), .ZN(
        n47) );
  AND2_X1 U18 ( .A1(warp_checker_fence_regs_wr_fence_en[21]), .A2(n225), .ZN(
        n48) );
  AND2_X1 U19 ( .A1(warp_checker_fence_regs_wr_fence_en[22]), .A2(n225), .ZN(
        n49) );
  AND2_X1 U20 ( .A1(warp_checker_fence_regs_wr_fence_en[23]), .A2(n223), .ZN(
        n50) );
  AND2_X1 U21 ( .A1(warp_checker_fence_regs_wr_fence_en[24]), .A2(n225), .ZN(
        n51) );
  AND2_X1 U22 ( .A1(warp_checker_fence_regs_wr_fence_en[25]), .A2(n223), .ZN(
        n52) );
  AND2_X1 U23 ( .A1(warp_checker_fence_regs_wr_fence_en[26]), .A2(n225), .ZN(
        n53) );
  AND2_X1 U24 ( .A1(warp_checker_fence_regs_wr_fence_en[27]), .A2(n225), .ZN(
        n54) );
  AND2_X1 U25 ( .A1(warp_checker_fence_regs_wr_fence_en[0]), .A2(n223), .ZN(
        n55) );
  AND2_X1 U26 ( .A1(warp_checker_fence_regs_wr_fence_en[3]), .A2(n224), .ZN(
        n56) );
  AND2_X1 U27 ( .A1(warp_checker_fence_regs_wr_fence_en[9]), .A2(n224), .ZN(
        n57) );
  AND2_X1 U28 ( .A1(warp_checker_fence_regs_wr_fence_en[15]), .A2(n224), .ZN(
        n58) );
  AND2_X1 U29 ( .A1(warp_checker_fence_regs_wr_fence_en[28]), .A2(n224), .ZN(
        n59) );
  AND2_X1 U30 ( .A1(warp_checker_fence_regs_wr_fence_en[29]), .A2(n224), .ZN(
        n60) );
  AND2_X1 U31 ( .A1(warp_checker_fence_regs_wr_fence_en[31]), .A2(n224), .ZN(
        n61) );
  AND2_X1 U32 ( .A1(warp_checker_fence_regs_wr_fence_en[12]), .A2(n226), .ZN(
        n62) );
  AND2_X1 U33 ( .A1(warp_checker_fence_regs_wr_fence_en[17]), .A2(n226), .ZN(
        n63) );
  AND2_X1 U34 ( .A1(warp_checker_fence_regs_wr_fence_en[30]), .A2(n226), .ZN(
        n64) );
  INV_X1 U35 ( .A(n220), .ZN(n164) );
  INV_X1 U36 ( .A(n219), .ZN(n175) );
  INV_X1 U37 ( .A(n219), .ZN(n163) );
  INV_X1 U38 ( .A(n218), .ZN(n160) );
  INV_X1 U39 ( .A(n219), .ZN(n172) );
  INV_X1 U40 ( .A(n220), .ZN(n170) );
  INV_X1 U41 ( .A(n220), .ZN(n171) );
  INV_X1 U42 ( .A(n219), .ZN(n174) );
  INV_X1 U43 ( .A(n218), .ZN(n165) );
  INV_X1 U44 ( .A(n218), .ZN(n167) );
  INV_X1 U45 ( .A(n221), .ZN(n178) );
  INV_X1 U46 ( .A(n221), .ZN(n177) );
  BUF_X1 U47 ( .A(n229), .Z(n218) );
  BUF_X1 U48 ( .A(n237), .Z(n189) );
  BUF_X1 U49 ( .A(n232), .Z(n204) );
  BUF_X1 U50 ( .A(n235), .Z(n196) );
  BUF_X1 U51 ( .A(n234), .Z(n197) );
  BUF_X1 U52 ( .A(n237), .Z(n190) );
  BUF_X1 U53 ( .A(n235), .Z(n194) );
  BUF_X1 U54 ( .A(n236), .Z(n193) );
  BUF_X1 U55 ( .A(n236), .Z(n192) );
  BUF_X1 U56 ( .A(n230), .Z(n210) );
  BUF_X1 U57 ( .A(n230), .Z(n217) );
  BUF_X1 U58 ( .A(n230), .Z(n216) );
  BUF_X1 U59 ( .A(n235), .Z(n195) );
  BUF_X1 U60 ( .A(n236), .Z(n191) );
  BUF_X1 U61 ( .A(n231), .Z(n209) );
  BUF_X1 U62 ( .A(n234), .Z(n199) );
  BUF_X1 U63 ( .A(n234), .Z(n198) );
  BUF_X1 U64 ( .A(n231), .Z(n207) );
  BUF_X1 U65 ( .A(n231), .Z(n206) );
  BUF_X1 U66 ( .A(n232), .Z(n205) );
  BUF_X1 U67 ( .A(n233), .Z(n202) );
  BUF_X1 U68 ( .A(n233), .Z(n201) );
  BUF_X1 U69 ( .A(n233), .Z(n200) );
  BUF_X1 U70 ( .A(n232), .Z(n203) );
  BUF_X1 U71 ( .A(n229), .Z(n220) );
  BUF_X1 U72 ( .A(n229), .Z(n219) );
  BUF_X1 U73 ( .A(n228), .Z(n221) );
  BUF_X1 U74 ( .A(n238), .Z(n186) );
  BUF_X1 U75 ( .A(n239), .Z(n183) );
  BUF_X1 U76 ( .A(n238), .Z(n187) );
  BUF_X1 U77 ( .A(n239), .Z(n182) );
  BUF_X1 U78 ( .A(n239), .Z(n184) );
  BUF_X1 U79 ( .A(n237), .Z(n188) );
  BUF_X1 U80 ( .A(n238), .Z(n185) );
  BUF_X1 U81 ( .A(n240), .Z(n181) );
  BUF_X1 U82 ( .A(n228), .Z(n222) );
  BUF_X1 U83 ( .A(n227), .Z(n225) );
  BUF_X1 U84 ( .A(n227), .Z(n224) );
  BUF_X1 U85 ( .A(n228), .Z(n223) );
  BUF_X1 U86 ( .A(n227), .Z(n226) );
  BUF_X1 U87 ( .A(n240), .Z(n179) );
  BUF_X1 U88 ( .A(n240), .Z(n180) );
  BUF_X1 U89 ( .A(n244), .Z(n234) );
  BUF_X1 U90 ( .A(n243), .Z(n235) );
  BUF_X1 U91 ( .A(n243), .Z(n236) );
  BUF_X1 U92 ( .A(n242), .Z(n237) );
  BUF_X1 U93 ( .A(n244), .Z(n233) );
  BUF_X1 U94 ( .A(n246), .Z(n230) );
  BUF_X1 U95 ( .A(n245), .Z(n231) );
  BUF_X1 U96 ( .A(n245), .Z(n232) );
  BUF_X1 U97 ( .A(n246), .Z(n229) );
  BUF_X1 U98 ( .A(n241), .Z(n239) );
  BUF_X1 U99 ( .A(n242), .Z(n238) );
  BUF_X1 U100 ( .A(n241), .Z(n240) );
  BUF_X1 U101 ( .A(n247), .Z(n227) );
  BUF_X1 U102 ( .A(n247), .Z(n228) );
  INV_X1 U103 ( .A(n158), .ZN(n244) );
  INV_X1 U104 ( .A(n158), .ZN(n243) );
  INV_X1 U105 ( .A(n158), .ZN(n242) );
  INV_X1 U106 ( .A(n159), .ZN(n246) );
  INV_X1 U107 ( .A(n159), .ZN(n245) );
  INV_X1 U108 ( .A(n158), .ZN(n241) );
  INV_X1 U109 ( .A(n159), .ZN(n247) );
  BUF_X1 U110 ( .A(warp_scheduler_reset), .Z(n158) );
  BUF_X1 U111 ( .A(warp_scheduler_reset), .Z(n159) );
  AND2_X1 U112 ( .A1(fence_regs_rd_fence_en[1]), .A2(n201), .ZN(
        warp_checker_fence_regs_rd_fence_en[1]) );
  AND2_X1 U113 ( .A1(fence_regs_rd_fence_en[0]), .A2(n199), .ZN(
        warp_checker_fence_regs_rd_fence_en[0]) );
  AND2_X1 U114 ( .A1(fence_regs_rd_fence_en[22]), .A2(n201), .ZN(
        warp_checker_fence_regs_rd_fence_en[22]) );
  AND2_X1 U115 ( .A1(fence_regs_rd_fence_en[18]), .A2(n201), .ZN(
        warp_checker_fence_regs_rd_fence_en[18]) );
  AND2_X1 U116 ( .A1(fence_regs_rd_fence_en[14]), .A2(n200), .ZN(
        warp_checker_fence_regs_rd_fence_en[14]) );
  AND2_X1 U117 ( .A1(fence_regs_rd_fence_en[9]), .A2(n189), .ZN(
        warp_checker_fence_regs_rd_fence_en[9]) );
  AND2_X1 U118 ( .A1(fence_regs_rd_fence_en[26]), .A2(n202), .ZN(
        warp_checker_fence_regs_rd_fence_en[26]) );
  AND2_X1 U119 ( .A1(fence_regs_rd_fence_en[30]), .A2(n203), .ZN(
        warp_checker_fence_regs_rd_fence_en[30]) );
  AND2_X1 U120 ( .A1(fence_regs_rd_fence_en[31]), .A2(n203), .ZN(
        warp_checker_fence_regs_rd_fence_en[31]) );
  AND2_X1 U121 ( .A1(fence_regs_rd_fence_en[2]), .A2(n203), .ZN(
        warp_checker_fence_regs_rd_fence_en[2]) );
  AND2_X1 U122 ( .A1(fence_regs_rd_fence_en[16]), .A2(n200), .ZN(
        warp_checker_fence_regs_rd_fence_en[16]) );
  AND2_X1 U123 ( .A1(fence_regs_rd_fence_en[15]), .A2(n200), .ZN(
        warp_checker_fence_regs_rd_fence_en[15]) );
  AND2_X1 U124 ( .A1(fence_regs_rd_fence_en[11]), .A2(n200), .ZN(
        warp_checker_fence_regs_rd_fence_en[11]) );
  AND2_X1 U125 ( .A1(fence_regs_rd_fence_en[23]), .A2(n202), .ZN(
        warp_checker_fence_regs_rd_fence_en[23]) );
  AND2_X1 U126 ( .A1(fence_regs_rd_fence_en[19]), .A2(n201), .ZN(
        warp_checker_fence_regs_rd_fence_en[19]) );
  AND2_X1 U127 ( .A1(fence_regs_rd_fence_en[29]), .A2(n202), .ZN(
        warp_checker_fence_regs_rd_fence_en[29]) );
  AND2_X1 U128 ( .A1(fence_regs_rd_fence_en[28]), .A2(n202), .ZN(
        warp_checker_fence_regs_rd_fence_en[28]) );
  AND2_X1 U129 ( .A1(fence_regs_rd_fence_en[27]), .A2(n202), .ZN(
        warp_checker_fence_regs_rd_fence_en[27]) );
  AND2_X1 U130 ( .A1(fence_regs_rd_fence_en[17]), .A2(n201), .ZN(
        warp_checker_fence_regs_rd_fence_en[17]) );
  AND2_X1 U131 ( .A1(fence_regs_rd_fence_en[7]), .A2(n204), .ZN(
        warp_checker_fence_regs_rd_fence_en[7]) );
  AND2_X1 U132 ( .A1(fence_regs_rd_fence_en[10]), .A2(n200), .ZN(
        warp_checker_fence_regs_rd_fence_en[10]) );
  AND2_X1 U133 ( .A1(fence_regs_rd_fence_en[13]), .A2(n200), .ZN(
        warp_checker_fence_regs_rd_fence_en[13]) );
  AND2_X1 U134 ( .A1(fence_regs_rd_fence_en[12]), .A2(n200), .ZN(
        warp_checker_fence_regs_rd_fence_en[12]) );
  AND2_X1 U135 ( .A1(fence_regs_rd_fence_en[25]), .A2(n202), .ZN(
        warp_checker_fence_regs_rd_fence_en[25]) );
  AND2_X1 U136 ( .A1(fence_regs_rd_fence_en[24]), .A2(n202), .ZN(
        warp_checker_fence_regs_rd_fence_en[24]) );
  AND2_X1 U137 ( .A1(fence_regs_rd_fence_en[21]), .A2(n201), .ZN(
        warp_checker_fence_regs_rd_fence_en[21]) );
  AND2_X1 U138 ( .A1(fence_regs_rd_fence_en[20]), .A2(n201), .ZN(
        warp_checker_fence_regs_rd_fence_en[20]) );
  AND2_X1 U139 ( .A1(fence_regs_rd_fence_en[8]), .A2(n204), .ZN(
        warp_checker_fence_regs_rd_fence_en[8]) );
  AND2_X1 U140 ( .A1(fence_regs_rd_fence_en[3]), .A2(n203), .ZN(
        warp_checker_fence_regs_rd_fence_en[3]) );
  AND2_X1 U141 ( .A1(fence_regs_rd_fence_en[4]), .A2(n203), .ZN(
        warp_checker_fence_regs_rd_fence_en[4]) );
  AND2_X1 U142 ( .A1(\fence_regs_rd_cta_id[21><2] ), .A2(n218), .ZN(
        \warp_checker_fence_regs_rd_cta_id[21><2] ) );
  AND2_X1 U143 ( .A1(fence_regs_rd_fence_en[5]), .A2(n203), .ZN(
        warp_checker_fence_regs_rd_fence_en[5]) );
  AND2_X1 U144 ( .A1(fence_regs_rd_fence_en[6]), .A2(n203), .ZN(
        warp_checker_fence_regs_rd_fence_en[6]) );
  AND2_X1 U145 ( .A1(\fence_regs_rd_cta_id[22><1] ), .A2(n218), .ZN(
        \warp_checker_fence_regs_rd_cta_id[22><1] ) );
  AND2_X1 U146 ( .A1(\fence_regs_rd_cta_id[22><0] ), .A2(n218), .ZN(
        \warp_checker_fence_regs_rd_cta_id[22><0] ) );
  AND2_X1 U147 ( .A1(\fence_regs_rd_cta_id[21><3] ), .A2(n218), .ZN(
        \warp_checker_fence_regs_rd_cta_id[21><3] ) );
  AND2_X1 U148 ( .A1(\fence_regs_rd_cta_id[23><1] ), .A2(n189), .ZN(
        \warp_checker_fence_regs_rd_cta_id[23><1] ) );
  AND2_X1 U149 ( .A1(\fence_regs_rd_cta_id[0><1] ), .A2(n204), .ZN(
        \warp_checker_fence_regs_rd_cta_id[0><1] ) );
  AND2_X1 U150 ( .A1(\fence_regs_rd_cta_id[0><2] ), .A2(n204), .ZN(
        \warp_checker_fence_regs_rd_cta_id[0><2] ) );
  AND2_X1 U151 ( .A1(\fence_regs_rd_cta_id[0><3] ), .A2(n204), .ZN(
        \warp_checker_fence_regs_rd_cta_id[0><3] ) );
  AND2_X1 U152 ( .A1(\fence_regs_rd_cta_id[5><1] ), .A2(n197), .ZN(
        \warp_checker_fence_regs_rd_cta_id[5><1] ) );
  AND2_X1 U153 ( .A1(\fence_regs_rd_cta_id[5><2] ), .A2(n197), .ZN(
        \warp_checker_fence_regs_rd_cta_id[5><2] ) );
  AND2_X1 U154 ( .A1(\fence_regs_rd_cta_id[5><3] ), .A2(n197), .ZN(
        \warp_checker_fence_regs_rd_cta_id[5><3] ) );
  AND2_X1 U155 ( .A1(\fence_regs_rd_cta_id[4><1] ), .A2(n196), .ZN(
        \warp_checker_fence_regs_rd_cta_id[4><1] ) );
  AND2_X1 U156 ( .A1(\fence_regs_rd_cta_id[4><2] ), .A2(n196), .ZN(
        \warp_checker_fence_regs_rd_cta_id[4><2] ) );
  AND2_X1 U157 ( .A1(\fence_regs_rd_cta_id[4><3] ), .A2(n196), .ZN(
        \warp_checker_fence_regs_rd_cta_id[4><3] ) );
  AND2_X1 U158 ( .A1(\fence_regs_rd_cta_id[9><1] ), .A2(n199), .ZN(
        \warp_checker_fence_regs_rd_cta_id[9><1] ) );
  AND2_X1 U159 ( .A1(\fence_regs_rd_cta_id[9><2] ), .A2(n199), .ZN(
        \warp_checker_fence_regs_rd_cta_id[9><2] ) );
  AND2_X1 U160 ( .A1(\fence_regs_rd_cta_id[9><3] ), .A2(n199), .ZN(
        \warp_checker_fence_regs_rd_cta_id[9><3] ) );
  AND2_X1 U161 ( .A1(\fence_regs_rd_cta_id[0><0] ), .A2(n204), .ZN(
        \warp_checker_fence_regs_rd_cta_id[0><0] ) );
  AND2_X1 U162 ( .A1(\fence_regs_rd_cta_id[5><0] ), .A2(n197), .ZN(
        \warp_checker_fence_regs_rd_cta_id[5><0] ) );
  AND2_X1 U163 ( .A1(\fence_regs_rd_cta_id[4><0] ), .A2(n196), .ZN(
        \warp_checker_fence_regs_rd_cta_id[4><0] ) );
  AND2_X1 U164 ( .A1(\fence_regs_rd_cta_id[9><0] ), .A2(n199), .ZN(
        \warp_checker_fence_regs_rd_cta_id[9><0] ) );
  AND2_X1 U165 ( .A1(\fence_regs_rd_cta_id[3><1] ), .A2(n193), .ZN(
        \warp_checker_fence_regs_rd_cta_id[3><1] ) );
  AND2_X1 U166 ( .A1(\fence_regs_rd_cta_id[3><2] ), .A2(n196), .ZN(
        \warp_checker_fence_regs_rd_cta_id[3><2] ) );
  AND2_X1 U167 ( .A1(\fence_regs_rd_cta_id[3><3] ), .A2(n196), .ZN(
        \warp_checker_fence_regs_rd_cta_id[3><3] ) );
  AND2_X1 U168 ( .A1(\fence_regs_rd_cta_id[6><1] ), .A2(n197), .ZN(
        \warp_checker_fence_regs_rd_cta_id[6><1] ) );
  AND2_X1 U169 ( .A1(\fence_regs_rd_cta_id[6><2] ), .A2(n197), .ZN(
        \warp_checker_fence_regs_rd_cta_id[6><2] ) );
  AND2_X1 U170 ( .A1(\fence_regs_rd_cta_id[6><3] ), .A2(n198), .ZN(
        \warp_checker_fence_regs_rd_cta_id[6><3] ) );
  AND2_X1 U171 ( .A1(\fence_regs_rd_cta_id[14><1] ), .A2(n207), .ZN(
        \warp_checker_fence_regs_rd_cta_id[14><1] ) );
  AND2_X1 U172 ( .A1(\fence_regs_rd_cta_id[14><2] ), .A2(n207), .ZN(
        \warp_checker_fence_regs_rd_cta_id[14><2] ) );
  AND2_X1 U173 ( .A1(\fence_regs_rd_cta_id[14><3] ), .A2(n207), .ZN(
        \warp_checker_fence_regs_rd_cta_id[14><3] ) );
  AND2_X1 U174 ( .A1(\fence_regs_rd_cta_id[26><1] ), .A2(n191), .ZN(
        \warp_checker_fence_regs_rd_cta_id[26><1] ) );
  AND2_X1 U175 ( .A1(\fence_regs_rd_cta_id[26><2] ), .A2(n191), .ZN(
        \warp_checker_fence_regs_rd_cta_id[26><2] ) );
  AND2_X1 U176 ( .A1(\fence_regs_rd_cta_id[26><3] ), .A2(n194), .ZN(
        \warp_checker_fence_regs_rd_cta_id[26><3] ) );
  AND2_X1 U177 ( .A1(\fence_regs_rd_cta_id[30><1] ), .A2(n192), .ZN(
        \warp_checker_fence_regs_rd_cta_id[30><1] ) );
  AND2_X1 U178 ( .A1(\fence_regs_rd_cta_id[30><2] ), .A2(n194), .ZN(
        \warp_checker_fence_regs_rd_cta_id[30><2] ) );
  AND2_X1 U179 ( .A1(\fence_regs_rd_cta_id[30><3] ), .A2(n193), .ZN(
        \warp_checker_fence_regs_rd_cta_id[30><3] ) );
  AND2_X1 U180 ( .A1(\fence_regs_rd_cta_id[22><2] ), .A2(n196), .ZN(
        \warp_checker_fence_regs_rd_cta_id[22><2] ) );
  AND2_X1 U181 ( .A1(\fence_regs_rd_cta_id[22><3] ), .A2(n192), .ZN(
        \warp_checker_fence_regs_rd_cta_id[22><3] ) );
  AND2_X1 U182 ( .A1(\fence_regs_rd_cta_id[18><1] ), .A2(n210), .ZN(
        \warp_checker_fence_regs_rd_cta_id[18><1] ) );
  AND2_X1 U183 ( .A1(\fence_regs_rd_cta_id[18><2] ), .A2(n210), .ZN(
        \warp_checker_fence_regs_rd_cta_id[18><2] ) );
  AND2_X1 U184 ( .A1(\fence_regs_rd_cta_id[18><3] ), .A2(n216), .ZN(
        \warp_checker_fence_regs_rd_cta_id[18><3] ) );
  AND2_X1 U185 ( .A1(\fence_regs_rd_cta_id[3><0] ), .A2(n195), .ZN(
        \warp_checker_fence_regs_rd_cta_id[3><0] ) );
  AND2_X1 U186 ( .A1(\fence_regs_rd_cta_id[6><0] ), .A2(n197), .ZN(
        \warp_checker_fence_regs_rd_cta_id[6><0] ) );
  AND2_X1 U187 ( .A1(\fence_regs_rd_cta_id[14><0] ), .A2(n207), .ZN(
        \warp_checker_fence_regs_rd_cta_id[14><0] ) );
  AND2_X1 U188 ( .A1(\fence_regs_rd_cta_id[26><0] ), .A2(n190), .ZN(
        \warp_checker_fence_regs_rd_cta_id[26><0] ) );
  AND2_X1 U189 ( .A1(\fence_regs_rd_cta_id[30><0] ), .A2(n192), .ZN(
        \warp_checker_fence_regs_rd_cta_id[30><0] ) );
  AND2_X1 U190 ( .A1(\fence_regs_rd_cta_id[18><0] ), .A2(n210), .ZN(
        \warp_checker_fence_regs_rd_cta_id[18><0] ) );
  AND2_X1 U191 ( .A1(\fence_regs_rd_cta_id[1><1] ), .A2(n216), .ZN(
        \warp_checker_fence_regs_rd_cta_id[1><1] ) );
  AND2_X1 U192 ( .A1(\fence_regs_rd_cta_id[1><2] ), .A2(n216), .ZN(
        \warp_checker_fence_regs_rd_cta_id[1><2] ) );
  AND2_X1 U193 ( .A1(\fence_regs_rd_cta_id[1><3] ), .A2(n217), .ZN(
        \warp_checker_fence_regs_rd_cta_id[1><3] ) );
  AND2_X1 U194 ( .A1(\fence_regs_rd_cta_id[25><1] ), .A2(n190), .ZN(
        \warp_checker_fence_regs_rd_cta_id[25><1] ) );
  AND2_X1 U195 ( .A1(\fence_regs_rd_cta_id[25><2] ), .A2(n190), .ZN(
        \warp_checker_fence_regs_rd_cta_id[25><2] ) );
  AND2_X1 U196 ( .A1(\fence_regs_rd_cta_id[25><3] ), .A2(n194), .ZN(
        \warp_checker_fence_regs_rd_cta_id[25><3] ) );
  AND2_X1 U197 ( .A1(\fence_regs_rd_cta_id[24><1] ), .A2(n193), .ZN(
        \warp_checker_fence_regs_rd_cta_id[24><1] ) );
  AND2_X1 U198 ( .A1(\fence_regs_rd_cta_id[24><2] ), .A2(n190), .ZN(
        \warp_checker_fence_regs_rd_cta_id[24><2] ) );
  AND2_X1 U199 ( .A1(\fence_regs_rd_cta_id[24><3] ), .A2(n190), .ZN(
        \warp_checker_fence_regs_rd_cta_id[24><3] ) );
  AND2_X1 U200 ( .A1(\fence_regs_rd_cta_id[23><2] ), .A2(n193), .ZN(
        \warp_checker_fence_regs_rd_cta_id[23><2] ) );
  AND2_X1 U201 ( .A1(\fence_regs_rd_cta_id[23><3] ), .A2(n190), .ZN(
        \warp_checker_fence_regs_rd_cta_id[23><3] ) );
  AND2_X1 U202 ( .A1(\fence_regs_rd_cta_id[21><0] ), .A2(n217), .ZN(
        \warp_checker_fence_regs_rd_cta_id[21><0] ) );
  AND2_X1 U203 ( .A1(\fence_regs_rd_cta_id[21><1] ), .A2(n217), .ZN(
        \warp_checker_fence_regs_rd_cta_id[21><1] ) );
  AND2_X1 U204 ( .A1(\fence_regs_rd_cta_id[20><1] ), .A2(n217), .ZN(
        \warp_checker_fence_regs_rd_cta_id[20><1] ) );
  AND2_X1 U205 ( .A1(\fence_regs_rd_cta_id[20><2] ), .A2(n217), .ZN(
        \warp_checker_fence_regs_rd_cta_id[20><2] ) );
  AND2_X1 U206 ( .A1(\fence_regs_rd_cta_id[20><3] ), .A2(n217), .ZN(
        \warp_checker_fence_regs_rd_cta_id[20><3] ) );
  AND2_X1 U207 ( .A1(\fence_regs_rd_cta_id[19><1] ), .A2(n209), .ZN(
        \warp_checker_fence_regs_rd_cta_id[19><1] ) );
  AND2_X1 U208 ( .A1(\fence_regs_rd_cta_id[19><2] ), .A2(n216), .ZN(
        \warp_checker_fence_regs_rd_cta_id[19><2] ) );
  AND2_X1 U209 ( .A1(\fence_regs_rd_cta_id[19><3] ), .A2(n216), .ZN(
        \warp_checker_fence_regs_rd_cta_id[19><3] ) );
  AND2_X1 U210 ( .A1(\fence_regs_rd_cta_id[29><1] ), .A2(n195), .ZN(
        \warp_checker_fence_regs_rd_cta_id[29><1] ) );
  AND2_X1 U211 ( .A1(\fence_regs_rd_cta_id[29><2] ), .A2(n192), .ZN(
        \warp_checker_fence_regs_rd_cta_id[29><2] ) );
  AND2_X1 U212 ( .A1(\fence_regs_rd_cta_id[29><3] ), .A2(n192), .ZN(
        \warp_checker_fence_regs_rd_cta_id[29><3] ) );
  AND2_X1 U213 ( .A1(\fence_regs_rd_cta_id[28><1] ), .A2(n191), .ZN(
        \warp_checker_fence_regs_rd_cta_id[28><1] ) );
  AND2_X1 U214 ( .A1(\fence_regs_rd_cta_id[28><2] ), .A2(n194), .ZN(
        \warp_checker_fence_regs_rd_cta_id[28><2] ) );
  AND2_X1 U215 ( .A1(\fence_regs_rd_cta_id[28><3] ), .A2(n195), .ZN(
        \warp_checker_fence_regs_rd_cta_id[28><3] ) );
  AND2_X1 U216 ( .A1(\fence_regs_rd_cta_id[27><1] ), .A2(n191), .ZN(
        \warp_checker_fence_regs_rd_cta_id[27><1] ) );
  AND2_X1 U217 ( .A1(\fence_regs_rd_cta_id[27><2] ), .A2(n191), .ZN(
        \warp_checker_fence_regs_rd_cta_id[27><2] ) );
  AND2_X1 U218 ( .A1(\fence_regs_rd_cta_id[27><3] ), .A2(n194), .ZN(
        \warp_checker_fence_regs_rd_cta_id[27><3] ) );
  AND2_X1 U219 ( .A1(\fence_regs_rd_cta_id[17><1] ), .A2(n210), .ZN(
        \warp_checker_fence_regs_rd_cta_id[17><1] ) );
  AND2_X1 U220 ( .A1(\fence_regs_rd_cta_id[17><2] ), .A2(n210), .ZN(
        \warp_checker_fence_regs_rd_cta_id[17><2] ) );
  AND2_X1 U221 ( .A1(\fence_regs_rd_cta_id[17><3] ), .A2(n210), .ZN(
        \warp_checker_fence_regs_rd_cta_id[17><3] ) );
  AND2_X1 U222 ( .A1(\fence_regs_rd_cta_id[16><1] ), .A2(n209), .ZN(
        \warp_checker_fence_regs_rd_cta_id[16><1] ) );
  AND2_X1 U223 ( .A1(\fence_regs_rd_cta_id[16><2] ), .A2(n209), .ZN(
        \warp_checker_fence_regs_rd_cta_id[16><2] ) );
  AND2_X1 U224 ( .A1(\fence_regs_rd_cta_id[16><3] ), .A2(n209), .ZN(
        \warp_checker_fence_regs_rd_cta_id[16><3] ) );
  AND2_X1 U225 ( .A1(\fence_regs_rd_cta_id[15><1] ), .A2(n207), .ZN(
        \warp_checker_fence_regs_rd_cta_id[15><1] ) );
  AND2_X1 U226 ( .A1(\fence_regs_rd_cta_id[15><2] ), .A2(n209), .ZN(
        \warp_checker_fence_regs_rd_cta_id[15><2] ) );
  AND2_X1 U227 ( .A1(\fence_regs_rd_cta_id[15><3] ), .A2(n209), .ZN(
        \warp_checker_fence_regs_rd_cta_id[15><3] ) );
  AND2_X1 U228 ( .A1(\fence_regs_rd_cta_id[10><1] ), .A2(n205), .ZN(
        \warp_checker_fence_regs_rd_cta_id[10><1] ) );
  AND2_X1 U229 ( .A1(\fence_regs_rd_cta_id[10><2] ), .A2(n205), .ZN(
        \warp_checker_fence_regs_rd_cta_id[10><2] ) );
  AND2_X1 U230 ( .A1(\fence_regs_rd_cta_id[10><3] ), .A2(n205), .ZN(
        \warp_checker_fence_regs_rd_cta_id[10><3] ) );
  AND2_X1 U231 ( .A1(\fence_regs_rd_cta_id[8><1] ), .A2(n198), .ZN(
        \warp_checker_fence_regs_rd_cta_id[8><1] ) );
  AND2_X1 U232 ( .A1(\fence_regs_rd_cta_id[8><2] ), .A2(n199), .ZN(
        \warp_checker_fence_regs_rd_cta_id[8><2] ) );
  AND2_X1 U233 ( .A1(\fence_regs_rd_cta_id[8><3] ), .A2(n199), .ZN(
        \warp_checker_fence_regs_rd_cta_id[8><3] ) );
  AND2_X1 U234 ( .A1(\fence_regs_rd_cta_id[7><1] ), .A2(n198), .ZN(
        \warp_checker_fence_regs_rd_cta_id[7><1] ) );
  AND2_X1 U235 ( .A1(\fence_regs_rd_cta_id[7><2] ), .A2(n198), .ZN(
        \warp_checker_fence_regs_rd_cta_id[7><2] ) );
  AND2_X1 U236 ( .A1(\fence_regs_rd_cta_id[7><3] ), .A2(n198), .ZN(
        \warp_checker_fence_regs_rd_cta_id[7><3] ) );
  AND2_X1 U237 ( .A1(\fence_regs_rd_cta_id[13><1] ), .A2(n206), .ZN(
        \warp_checker_fence_regs_rd_cta_id[13><1] ) );
  AND2_X1 U238 ( .A1(\fence_regs_rd_cta_id[13><2] ), .A2(n206), .ZN(
        \warp_checker_fence_regs_rd_cta_id[13><2] ) );
  AND2_X1 U239 ( .A1(\fence_regs_rd_cta_id[13><3] ), .A2(n207), .ZN(
        \warp_checker_fence_regs_rd_cta_id[13><3] ) );
  AND2_X1 U240 ( .A1(\fence_regs_rd_cta_id[12><1] ), .A2(n206), .ZN(
        \warp_checker_fence_regs_rd_cta_id[12><1] ) );
  AND2_X1 U241 ( .A1(\fence_regs_rd_cta_id[12><2] ), .A2(n206), .ZN(
        \warp_checker_fence_regs_rd_cta_id[12><2] ) );
  AND2_X1 U242 ( .A1(\fence_regs_rd_cta_id[12><3] ), .A2(n206), .ZN(
        \warp_checker_fence_regs_rd_cta_id[12><3] ) );
  AND2_X1 U243 ( .A1(\fence_regs_rd_cta_id[11><1] ), .A2(n205), .ZN(
        \warp_checker_fence_regs_rd_cta_id[11><1] ) );
  AND2_X1 U244 ( .A1(\fence_regs_rd_cta_id[11><2] ), .A2(n205), .ZN(
        \warp_checker_fence_regs_rd_cta_id[11><2] ) );
  AND2_X1 U245 ( .A1(\fence_regs_rd_cta_id[11><3] ), .A2(n205), .ZN(
        \warp_checker_fence_regs_rd_cta_id[11><3] ) );
  AND2_X1 U246 ( .A1(\fence_regs_rd_cta_id[1><0] ), .A2(n216), .ZN(
        \warp_checker_fence_regs_rd_cta_id[1><0] ) );
  AND2_X1 U247 ( .A1(\fence_regs_rd_cta_id[2><1] ), .A2(n192), .ZN(
        \warp_checker_fence_regs_rd_cta_id[2><1] ) );
  AND2_X1 U248 ( .A1(\fence_regs_rd_cta_id[2><2] ), .A2(n192), .ZN(
        \warp_checker_fence_regs_rd_cta_id[2><2] ) );
  AND2_X1 U249 ( .A1(\fence_regs_rd_cta_id[2><3] ), .A2(n195), .ZN(
        \warp_checker_fence_regs_rd_cta_id[2><3] ) );
  AND2_X1 U250 ( .A1(\fence_regs_rd_cta_id[31><1] ), .A2(n195), .ZN(
        \warp_checker_fence_regs_rd_cta_id[31><1] ) );
  AND2_X1 U251 ( .A1(\fence_regs_rd_cta_id[31><2] ), .A2(n193), .ZN(
        \warp_checker_fence_regs_rd_cta_id[31><2] ) );
  AND2_X1 U252 ( .A1(\fence_regs_rd_cta_id[31><3] ), .A2(n195), .ZN(
        \warp_checker_fence_regs_rd_cta_id[31><3] ) );
  AND2_X1 U253 ( .A1(\fence_regs_rd_cta_id[25><0] ), .A2(n195), .ZN(
        \warp_checker_fence_regs_rd_cta_id[25><0] ) );
  AND2_X1 U254 ( .A1(\fence_regs_rd_cta_id[24><0] ), .A2(n190), .ZN(
        \warp_checker_fence_regs_rd_cta_id[24><0] ) );
  AND2_X1 U255 ( .A1(\fence_regs_rd_cta_id[23><0] ), .A2(n193), .ZN(
        \warp_checker_fence_regs_rd_cta_id[23><0] ) );
  AND2_X1 U256 ( .A1(\fence_regs_rd_cta_id[20><0] ), .A2(n217), .ZN(
        \warp_checker_fence_regs_rd_cta_id[20><0] ) );
  AND2_X1 U257 ( .A1(\fence_regs_rd_cta_id[19><0] ), .A2(n216), .ZN(
        \warp_checker_fence_regs_rd_cta_id[19><0] ) );
  AND2_X1 U258 ( .A1(\fence_regs_rd_cta_id[29><0] ), .A2(n191), .ZN(
        \warp_checker_fence_regs_rd_cta_id[29><0] ) );
  AND2_X1 U259 ( .A1(\fence_regs_rd_cta_id[28><0] ), .A2(n191), .ZN(
        \warp_checker_fence_regs_rd_cta_id[28><0] ) );
  AND2_X1 U260 ( .A1(\fence_regs_rd_cta_id[27><0] ), .A2(n194), .ZN(
        \warp_checker_fence_regs_rd_cta_id[27><0] ) );
  AND2_X1 U261 ( .A1(\fence_regs_rd_cta_id[17><0] ), .A2(n210), .ZN(
        \warp_checker_fence_regs_rd_cta_id[17><0] ) );
  AND2_X1 U262 ( .A1(\fence_regs_rd_cta_id[16><0] ), .A2(n209), .ZN(
        \warp_checker_fence_regs_rd_cta_id[16><0] ) );
  AND2_X1 U263 ( .A1(\fence_regs_rd_cta_id[15><0] ), .A2(n207), .ZN(
        \warp_checker_fence_regs_rd_cta_id[15><0] ) );
  AND2_X1 U264 ( .A1(\fence_regs_rd_cta_id[10><0] ), .A2(n204), .ZN(
        \warp_checker_fence_regs_rd_cta_id[10><0] ) );
  AND2_X1 U265 ( .A1(\fence_regs_rd_cta_id[8><0] ), .A2(n198), .ZN(
        \warp_checker_fence_regs_rd_cta_id[8><0] ) );
  AND2_X1 U266 ( .A1(\fence_regs_rd_cta_id[7><0] ), .A2(n198), .ZN(
        \warp_checker_fence_regs_rd_cta_id[7><0] ) );
  AND2_X1 U267 ( .A1(\fence_regs_rd_cta_id[13><0] ), .A2(n206), .ZN(
        \warp_checker_fence_regs_rd_cta_id[13><0] ) );
  AND2_X1 U268 ( .A1(\fence_regs_rd_cta_id[12><0] ), .A2(n206), .ZN(
        \warp_checker_fence_regs_rd_cta_id[12><0] ) );
  AND2_X1 U269 ( .A1(\fence_regs_rd_cta_id[11><0] ), .A2(n205), .ZN(
        \warp_checker_fence_regs_rd_cta_id[11><0] ) );
  AND2_X1 U270 ( .A1(\fence_regs_rd_cta_id[2><0] ), .A2(n194), .ZN(
        \warp_checker_fence_regs_rd_cta_id[2><0] ) );
  AND2_X1 U271 ( .A1(\fence_regs_rd_cta_id[31><0] ), .A2(n193), .ZN(
        \warp_checker_fence_regs_rd_cta_id[31><0] ) );
  AND2_X1 U272 ( .A1(warp_gen_fence_regs_cta_id_ld[3]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[3]) );
  AND2_X1 U273 ( .A1(warp_gen_fence_regs_cta_id_ld[4]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[4]) );
  AND2_X1 U274 ( .A1(warp_gen_fence_regs_cta_id_ld[5]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[5]) );
  AND2_X1 U275 ( .A1(warp_gen_fence_regs_cta_id_ld[6]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[6]) );
  AND2_X1 U276 ( .A1(warp_gen_fence_regs_cta_id_ld[7]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[7]) );
  AND2_X1 U277 ( .A1(warp_gen_fence_regs_cta_id_ld[8]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[8]) );
  AND2_X1 U278 ( .A1(warp_gen_fence_regs_cta_id_ld[9]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[9]) );
  AND2_X1 U279 ( .A1(warp_gen_fence_regs_cta_id_ld[30]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[30]) );
  AND2_X1 U280 ( .A1(warp_gen_fence_regs_cta_id_ld[31]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[31]) );
  AND2_X1 U281 ( .A1(warp_gen_fence_regs_cta_id_ld[10]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[10]) );
  AND2_X1 U282 ( .A1(warp_gen_fence_regs_cta_id_ld[11]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[11]) );
  AND2_X1 U283 ( .A1(warp_gen_fence_regs_cta_id_ld[12]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[12]) );
  AND2_X1 U284 ( .A1(warp_gen_fence_regs_cta_id_ld[13]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[13]) );
  AND2_X1 U285 ( .A1(warp_gen_fence_regs_cta_id_ld[14]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[14]) );
  AND2_X1 U286 ( .A1(warp_gen_fence_regs_cta_id_ld[15]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[15]) );
  AND2_X1 U287 ( .A1(warp_gen_fence_regs_cta_id_ld[16]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[16]) );
  AND2_X1 U288 ( .A1(warp_gen_fence_regs_cta_id_ld[0]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[0]) );
  AND2_X1 U289 ( .A1(warp_gen_fence_regs_cta_id_ld[1]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[1]) );
  AND2_X1 U290 ( .A1(warp_gen_fence_regs_cta_id_ld[2]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[2]) );
  AND2_X1 U291 ( .A1(warp_gen_fence_regs_cta_id_ld[17]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[17]) );
  AND2_X1 U292 ( .A1(warp_gen_fence_regs_cta_id_ld[18]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[18]) );
  AND2_X1 U293 ( .A1(warp_gen_fence_regs_cta_id_ld[19]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[19]) );
  AND2_X1 U294 ( .A1(warp_gen_fence_regs_cta_id_ld[20]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[20]) );
  AND2_X1 U295 ( .A1(warp_gen_fence_regs_cta_id_ld[21]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[21]) );
  AND2_X1 U296 ( .A1(warp_gen_fence_regs_cta_id_ld[22]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[22]) );
  AND2_X1 U297 ( .A1(warp_gen_fence_regs_cta_id_ld[23]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[23]) );
  AND2_X1 U298 ( .A1(warp_gen_fence_regs_cta_id_ld[24]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[24]) );
  AND2_X1 U299 ( .A1(warp_gen_fence_regs_cta_id_ld[25]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[25]) );
  AND2_X1 U300 ( .A1(warp_gen_fence_regs_cta_id_ld[26]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[26]) );
  AND2_X1 U301 ( .A1(warp_gen_fence_regs_cta_id_ld[27]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[27]) );
  AND2_X1 U302 ( .A1(warp_gen_fence_regs_cta_id_ld[28]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[28]) );
  AND2_X1 U303 ( .A1(warp_gen_fence_regs_cta_id_ld[29]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[29]) );
  AOI22_X1 U304 ( .A1(warp_checker_fence_regs_fence_en_ld[1]), .A2(n186), .B1(
        warp_gen_fence_regs_fence_en_ld[1]), .B2(n161), .ZN(n402) );
  AOI22_X1 U305 ( .A1(warp_checker_fence_regs_fence_en_ld[2]), .A2(n184), .B1(
        warp_gen_fence_regs_fence_en_ld[2]), .B2(n162), .ZN(n391) );
  AOI22_X1 U306 ( .A1(warp_checker_fence_regs_fence_en_ld[3]), .A2(n184), .B1(
        warp_gen_fence_regs_fence_en_ld[3]), .B2(n161), .ZN(n388) );
  AOI22_X1 U307 ( .A1(warp_checker_fence_regs_fence_en_ld[5]), .A2(n189), .B1(
        warp_gen_fence_regs_fence_en_ld[5]), .B2(n161), .ZN(n386) );
  AOI22_X1 U308 ( .A1(warp_checker_fence_regs_fence_en_ld[6]), .A2(n184), .B1(
        warp_gen_fence_regs_fence_en_ld[6]), .B2(n161), .ZN(n385) );
  AOI22_X1 U309 ( .A1(warp_checker_fence_regs_fence_en_ld[8]), .A2(n189), .B1(
        warp_gen_fence_regs_fence_en_ld[8]), .B2(n161), .ZN(n383) );
  AOI22_X1 U310 ( .A1(warp_checker_fence_regs_fence_en_ld[16]), .A2(n183), 
        .B1(warp_gen_fence_regs_fence_en_ld[16]), .B2(n162), .ZN(n406) );
  AOI22_X1 U311 ( .A1(warp_checker_fence_regs_fence_en_ld[17]), .A2(n186), 
        .B1(warp_gen_fence_regs_fence_en_ld[17]), .B2(n161), .ZN(n405) );
  AOI22_X1 U312 ( .A1(warp_checker_fence_regs_fence_en_ld[18]), .A2(n186), 
        .B1(warp_gen_fence_regs_fence_en_ld[18]), .B2(n162), .ZN(n404) );
  AOI22_X1 U313 ( .A1(warp_checker_fence_regs_fence_en_ld[19]), .A2(n183), 
        .B1(warp_gen_fence_regs_fence_en_ld[19]), .B2(n162), .ZN(n403) );
  AOI22_X1 U314 ( .A1(warp_checker_fence_regs_fence_en_ld[21]), .A2(n183), 
        .B1(warp_gen_fence_regs_fence_en_ld[21]), .B2(n162), .ZN(n400) );
  AOI22_X1 U315 ( .A1(warp_checker_fence_regs_fence_en_ld[22]), .A2(n187), 
        .B1(warp_gen_fence_regs_fence_en_ld[22]), .B2(n161), .ZN(n399) );
  AOI22_X1 U316 ( .A1(warp_checker_fence_regs_fence_en_ld[23]), .A2(n187), 
        .B1(warp_gen_fence_regs_fence_en_ld[23]), .B2(n162), .ZN(n398) );
  AOI22_X1 U317 ( .A1(warp_checker_fence_regs_fence_en_ld[24]), .A2(n183), 
        .B1(warp_gen_fence_regs_fence_en_ld[24]), .B2(n162), .ZN(n397) );
  AOI22_X1 U318 ( .A1(warp_checker_fence_regs_fence_en_ld[25]), .A2(n187), 
        .B1(warp_gen_fence_regs_fence_en_ld[25]), .B2(n161), .ZN(n396) );
  AOI22_X1 U319 ( .A1(warp_checker_fence_regs_fence_en_ld[26]), .A2(n188), 
        .B1(warp_gen_fence_regs_fence_en_ld[26]), .B2(n162), .ZN(n395) );
  AOI22_X1 U320 ( .A1(warp_checker_fence_regs_fence_en_ld[29]), .A2(n184), 
        .B1(warp_gen_fence_regs_fence_en_ld[29]), .B2(n162), .ZN(n392) );
  AOI22_X1 U321 ( .A1(warp_checker_fence_regs_fence_en_ld[31]), .A2(n188), 
        .B1(warp_gen_fence_regs_fence_en_ld[31]), .B2(n161), .ZN(n389) );
  AOI22_X1 U322 ( .A1(warp_checker_fence_regs_fence_en_ld[4]), .A2(n189), .B1(
        warp_gen_fence_regs_fence_en_ld[4]), .B2(n160), .ZN(n387) );
  AOI22_X1 U323 ( .A1(warp_checker_fence_regs_fence_en_ld[7]), .A2(n182), .B1(
        warp_gen_fence_regs_fence_en_ld[7]), .B2(n160), .ZN(n384) );
  AOI22_X1 U324 ( .A1(warp_checker_fence_regs_fence_en_ld[9]), .A2(n185), .B1(
        warp_gen_fence_regs_fence_en_ld[9]), .B2(n160), .ZN(n382) );
  AOI22_X1 U325 ( .A1(warp_checker_fence_regs_fence_en_ld[11]), .A2(n185), 
        .B1(warp_gen_fence_regs_fence_en_ld[11]), .B2(n160), .ZN(n411) );
  AOI22_X1 U326 ( .A1(warp_checker_fence_regs_fence_en_ld[14]), .A2(n182), 
        .B1(warp_gen_fence_regs_fence_en_ld[14]), .B2(n160), .ZN(n408) );
  AOI22_X1 U327 ( .A1(warp_checker_fence_regs_fence_en_ld[20]), .A2(n187), 
        .B1(warp_gen_fence_regs_fence_en_ld[20]), .B2(n160), .ZN(n401) );
  AOI22_X1 U328 ( .A1(warp_checker_fence_regs_fence_en_ld[27]), .A2(n182), 
        .B1(warp_gen_fence_regs_fence_en_ld[27]), .B2(n160), .ZN(n394) );
  AOI22_X1 U329 ( .A1(warp_checker_fence_regs_fence_en_ld[28]), .A2(n188), 
        .B1(warp_gen_fence_regs_fence_en_ld[28]), .B2(n160), .ZN(n393) );
  AOI22_X1 U330 ( .A1(warp_checker_fence_regs_fence_en_ld[30]), .A2(n188), 
        .B1(warp_gen_fence_regs_fence_en_ld[30]), .B2(n160), .ZN(n390) );
  AOI22_X1 U331 ( .A1(warp_checker_fence_regs_fence_en_ld[10]), .A2(n181), 
        .B1(warp_gen_fence_regs_fence_en_ld[10]), .B2(n163), .ZN(n412) );
  AOI22_X1 U332 ( .A1(warp_checker_fence_regs_fence_en_ld[12]), .A2(n185), 
        .B1(warp_gen_fence_regs_fence_en_ld[12]), .B2(n163), .ZN(n410) );
  AOI22_X1 U333 ( .A1(warp_checker_fence_regs_fence_en_ld[13]), .A2(n182), 
        .B1(warp_gen_fence_regs_fence_en_ld[13]), .B2(n163), .ZN(n409) );
  AOI22_X1 U334 ( .A1(warp_checker_fence_regs_fence_en_ld[15]), .A2(n186), 
        .B1(warp_gen_fence_regs_fence_en_ld[15]), .B2(n163), .ZN(n407) );
  AOI22_X1 U335 ( .A1(warp_checker_fence_regs_fence_en_ld[0]), .A2(n185), .B1(
        warp_gen_fence_regs_fence_en_ld[0]), .B2(n163), .ZN(n413) );
  AND2_X1 U336 ( .A1(\warp_gen_fence_regs_wr_cta_id[10><0] ), .A2(n173), .ZN(
        \fence_regs_wr_cta_id[10><0] ) );
  AND2_X1 U337 ( .A1(\warp_gen_fence_regs_wr_cta_id[11><0] ), .A2(n164), .ZN(
        \fence_regs_wr_cta_id[11><0] ) );
  AND2_X1 U338 ( .A1(\warp_gen_fence_regs_wr_cta_id[12><0] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[12><0] ) );
  AND2_X1 U339 ( .A1(\warp_gen_fence_regs_wr_cta_id[13><0] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[13><0] ) );
  AND2_X1 U340 ( .A1(\warp_gen_fence_regs_wr_cta_id[14><0] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[14><0] ) );
  AND2_X1 U341 ( .A1(\warp_gen_fence_regs_wr_cta_id[15><0] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[15><0] ) );
  AND2_X1 U342 ( .A1(\warp_gen_fence_regs_wr_cta_id[16><0] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[16><0] ) );
  AND2_X1 U343 ( .A1(\warp_gen_fence_regs_wr_cta_id[0><0] ), .A2(n173), .ZN(
        \fence_regs_wr_cta_id[0><0] ) );
  AND2_X1 U344 ( .A1(\warp_gen_fence_regs_wr_cta_id[1><0] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[1><0] ) );
  AND2_X1 U345 ( .A1(\warp_gen_fence_regs_wr_cta_id[2><0] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[2><0] ) );
  AND2_X1 U346 ( .A1(\warp_gen_fence_regs_wr_cta_id[17><0] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[17><0] ) );
  AND2_X1 U347 ( .A1(\warp_gen_fence_regs_wr_cta_id[18><0] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[18><0] ) );
  AND2_X1 U348 ( .A1(\warp_gen_fence_regs_wr_cta_id[19><0] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[19><0] ) );
  AND2_X1 U349 ( .A1(\warp_gen_fence_regs_wr_cta_id[20><0] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[20><0] ) );
  AND2_X1 U350 ( .A1(\warp_gen_fence_regs_wr_cta_id[21><0] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[21><0] ) );
  AND2_X1 U351 ( .A1(\warp_gen_fence_regs_wr_cta_id[22><0] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[22><0] ) );
  AND2_X1 U352 ( .A1(\warp_gen_fence_regs_wr_cta_id[23><0] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[23><0] ) );
  AND2_X1 U353 ( .A1(\warp_gen_fence_regs_wr_cta_id[24><0] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[24><0] ) );
  AND2_X1 U354 ( .A1(\warp_gen_fence_regs_wr_cta_id[25><0] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[25><0] ) );
  AND2_X1 U355 ( .A1(\warp_gen_fence_regs_wr_cta_id[26><0] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[26><0] ) );
  AND2_X1 U356 ( .A1(\warp_gen_fence_regs_wr_cta_id[27><0] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[27><0] ) );
  AND2_X1 U357 ( .A1(\warp_gen_fence_regs_wr_cta_id[28><0] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[28><0] ) );
  AND2_X1 U358 ( .A1(\warp_gen_fence_regs_wr_cta_id[29><0] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[29><0] ) );
  AND2_X1 U359 ( .A1(\warp_gen_fence_regs_wr_cta_id[10><1] ), .A2(n173), .ZN(
        \fence_regs_wr_cta_id[10><1] ) );
  AND2_X1 U360 ( .A1(\warp_gen_fence_regs_wr_cta_id[10><2] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[10><2] ) );
  AND2_X1 U361 ( .A1(\warp_gen_fence_regs_wr_cta_id[10><3] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[10><3] ) );
  AND2_X1 U362 ( .A1(\warp_gen_fence_regs_wr_cta_id[11><1] ), .A2(n164), .ZN(
        \fence_regs_wr_cta_id[11><1] ) );
  AND2_X1 U363 ( .A1(\warp_gen_fence_regs_wr_cta_id[11><2] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[11><2] ) );
  AND2_X1 U364 ( .A1(\warp_gen_fence_regs_wr_cta_id[11><3] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[11><3] ) );
  AND2_X1 U365 ( .A1(\warp_gen_fence_regs_wr_cta_id[12><1] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[12><1] ) );
  AND2_X1 U366 ( .A1(\warp_gen_fence_regs_wr_cta_id[12><2] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[12><2] ) );
  AND2_X1 U367 ( .A1(\warp_gen_fence_regs_wr_cta_id[12><3] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[12><3] ) );
  AND2_X1 U368 ( .A1(\warp_gen_fence_regs_wr_cta_id[13><1] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[13><1] ) );
  AND2_X1 U369 ( .A1(\warp_gen_fence_regs_wr_cta_id[13><2] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[13><2] ) );
  AND2_X1 U370 ( .A1(\warp_gen_fence_regs_wr_cta_id[13><3] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[13><3] ) );
  AND2_X1 U371 ( .A1(\warp_gen_fence_regs_wr_cta_id[14><1] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[14><1] ) );
  AND2_X1 U372 ( .A1(\warp_gen_fence_regs_wr_cta_id[14><2] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[14><2] ) );
  AND2_X1 U373 ( .A1(\warp_gen_fence_regs_wr_cta_id[14><3] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[14><3] ) );
  AND2_X1 U374 ( .A1(\warp_gen_fence_regs_wr_cta_id[15><1] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[15><1] ) );
  AND2_X1 U375 ( .A1(\warp_gen_fence_regs_wr_cta_id[15><2] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[15><2] ) );
  AND2_X1 U376 ( .A1(\warp_gen_fence_regs_wr_cta_id[15><3] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[15><3] ) );
  AND2_X1 U377 ( .A1(\warp_gen_fence_regs_wr_cta_id[16><1] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[16><1] ) );
  AND2_X1 U378 ( .A1(\warp_gen_fence_regs_wr_cta_id[16><2] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[16><2] ) );
  AND2_X1 U379 ( .A1(\warp_gen_fence_regs_wr_cta_id[16><3] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[16><3] ) );
  AND2_X1 U380 ( .A1(\warp_gen_fence_regs_wr_cta_id[0><1] ), .A2(n173), .ZN(
        \fence_regs_wr_cta_id[0><1] ) );
  AND2_X1 U381 ( .A1(\warp_gen_fence_regs_wr_cta_id[0><2] ), .A2(n173), .ZN(
        \fence_regs_wr_cta_id[0><2] ) );
  AND2_X1 U382 ( .A1(\warp_gen_fence_regs_wr_cta_id[0><3] ), .A2(n173), .ZN(
        \fence_regs_wr_cta_id[0><3] ) );
  AND2_X1 U383 ( .A1(\warp_gen_fence_regs_wr_cta_id[1><1] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[1><1] ) );
  AND2_X1 U384 ( .A1(\warp_gen_fence_regs_wr_cta_id[1><2] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[1><2] ) );
  AND2_X1 U385 ( .A1(\warp_gen_fence_regs_wr_cta_id[1><3] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[1><3] ) );
  AND2_X1 U386 ( .A1(\warp_gen_fence_regs_wr_cta_id[2><1] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[2><1] ) );
  AND2_X1 U387 ( .A1(\warp_gen_fence_regs_wr_cta_id[2><2] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[2><2] ) );
  AND2_X1 U388 ( .A1(\warp_gen_fence_regs_wr_cta_id[2><3] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[2><3] ) );
  AND2_X1 U389 ( .A1(\warp_gen_fence_regs_wr_cta_id[17><1] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[17><1] ) );
  AND2_X1 U390 ( .A1(\warp_gen_fence_regs_wr_cta_id[17><2] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[17><2] ) );
  AND2_X1 U391 ( .A1(\warp_gen_fence_regs_wr_cta_id[17><3] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[17><3] ) );
  AND2_X1 U392 ( .A1(\warp_gen_fence_regs_wr_cta_id[18><1] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[18><1] ) );
  AND2_X1 U393 ( .A1(\warp_gen_fence_regs_wr_cta_id[18><2] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[18><2] ) );
  AND2_X1 U394 ( .A1(\warp_gen_fence_regs_wr_cta_id[18><3] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[18><3] ) );
  AND2_X1 U395 ( .A1(\warp_gen_fence_regs_wr_cta_id[19><1] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[19><1] ) );
  AND2_X1 U396 ( .A1(\warp_gen_fence_regs_wr_cta_id[19><2] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[19><2] ) );
  AND2_X1 U397 ( .A1(\warp_gen_fence_regs_wr_cta_id[19><3] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[19><3] ) );
  AND2_X1 U398 ( .A1(\warp_gen_fence_regs_wr_cta_id[20><1] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[20><1] ) );
  AND2_X1 U399 ( .A1(\warp_gen_fence_regs_wr_cta_id[20><2] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[20><2] ) );
  AND2_X1 U400 ( .A1(\warp_gen_fence_regs_wr_cta_id[20><3] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[20><3] ) );
  AND2_X1 U401 ( .A1(\warp_gen_fence_regs_wr_cta_id[21><1] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[21><1] ) );
  AND2_X1 U402 ( .A1(\warp_gen_fence_regs_wr_cta_id[21><2] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[21><2] ) );
  AND2_X1 U403 ( .A1(\warp_gen_fence_regs_wr_cta_id[21><3] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[21><3] ) );
  AND2_X1 U404 ( .A1(\warp_gen_fence_regs_wr_cta_id[22><1] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[22><1] ) );
  AND2_X1 U405 ( .A1(\warp_gen_fence_regs_wr_cta_id[22><2] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[22><2] ) );
  AND2_X1 U406 ( .A1(\warp_gen_fence_regs_wr_cta_id[22><3] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[22><3] ) );
  AND2_X1 U407 ( .A1(\warp_gen_fence_regs_wr_cta_id[23><1] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[23><1] ) );
  AND2_X1 U408 ( .A1(\warp_gen_fence_regs_wr_cta_id[23><2] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[23><2] ) );
  AND2_X1 U409 ( .A1(\warp_gen_fence_regs_wr_cta_id[23><3] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[23><3] ) );
  AND2_X1 U410 ( .A1(\warp_gen_fence_regs_wr_cta_id[24><1] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[24><1] ) );
  AND2_X1 U411 ( .A1(\warp_gen_fence_regs_wr_cta_id[24><2] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[24><2] ) );
  AND2_X1 U412 ( .A1(\warp_gen_fence_regs_wr_cta_id[24><3] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[24><3] ) );
  AND2_X1 U413 ( .A1(\warp_gen_fence_regs_wr_cta_id[25><1] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[25><1] ) );
  AND2_X1 U414 ( .A1(\warp_gen_fence_regs_wr_cta_id[25><2] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[25><2] ) );
  AND2_X1 U415 ( .A1(\warp_gen_fence_regs_wr_cta_id[25><3] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[25><3] ) );
  AND2_X1 U416 ( .A1(\warp_gen_fence_regs_wr_cta_id[26><1] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[26><1] ) );
  AND2_X1 U417 ( .A1(\warp_gen_fence_regs_wr_cta_id[26><2] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[26><2] ) );
  AND2_X1 U418 ( .A1(\warp_gen_fence_regs_wr_cta_id[26><3] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[26><3] ) );
  AND2_X1 U419 ( .A1(\warp_gen_fence_regs_wr_cta_id[27><1] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[27><1] ) );
  AND2_X1 U420 ( .A1(\warp_gen_fence_regs_wr_cta_id[27><2] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[27><2] ) );
  AND2_X1 U421 ( .A1(\warp_gen_fence_regs_wr_cta_id[27><3] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[27><3] ) );
  AND2_X1 U422 ( .A1(\warp_gen_fence_regs_wr_cta_id[28><1] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[28><1] ) );
  AND2_X1 U423 ( .A1(\warp_gen_fence_regs_wr_cta_id[28><2] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[28><2] ) );
  AND2_X1 U424 ( .A1(\warp_gen_fence_regs_wr_cta_id[28><3] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[28><3] ) );
  AND2_X1 U425 ( .A1(\warp_gen_fence_regs_wr_cta_id[29><1] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[29><1] ) );
  AND2_X1 U426 ( .A1(\warp_gen_fence_regs_wr_cta_id[29><2] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[29><2] ) );
  AND2_X1 U427 ( .A1(\warp_gen_fence_regs_wr_cta_id[29><3] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[29><3] ) );
  INV_X1 U428 ( .A(n387), .ZN(n5) );
  INV_X1 U429 ( .A(n384), .ZN(n8) );
  INV_X1 U430 ( .A(n382), .ZN(n10) );
  INV_X1 U431 ( .A(n411), .ZN(n12) );
  INV_X1 U432 ( .A(n408), .ZN(n15) );
  INV_X1 U433 ( .A(n401), .ZN(n21) );
  INV_X1 U434 ( .A(n394), .ZN(n28) );
  INV_X1 U435 ( .A(n393), .ZN(n29) );
  INV_X1 U436 ( .A(n390), .ZN(n31) );
  AND2_X1 U437 ( .A1(\warp_gen_fence_regs_wr_cta_id[3><0] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[3><0] ) );
  AND2_X1 U438 ( .A1(\warp_gen_fence_regs_wr_cta_id[3><1] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[3><1] ) );
  AND2_X1 U439 ( .A1(\warp_gen_fence_regs_wr_cta_id[3><2] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[3><2] ) );
  AND2_X1 U440 ( .A1(\warp_gen_fence_regs_wr_cta_id[3><3] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[3><3] ) );
  AND2_X1 U441 ( .A1(\warp_gen_fence_regs_wr_cta_id[4><0] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[4><0] ) );
  AND2_X1 U442 ( .A1(\warp_gen_fence_regs_wr_cta_id[4><1] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[4><1] ) );
  AND2_X1 U443 ( .A1(\warp_gen_fence_regs_wr_cta_id[4><2] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[4><2] ) );
  AND2_X1 U444 ( .A1(\warp_gen_fence_regs_wr_cta_id[4><3] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[4><3] ) );
  AND2_X1 U445 ( .A1(\warp_gen_fence_regs_wr_cta_id[5><0] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[5><0] ) );
  AND2_X1 U446 ( .A1(\warp_gen_fence_regs_wr_cta_id[5><1] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[5><1] ) );
  AND2_X1 U447 ( .A1(\warp_gen_fence_regs_wr_cta_id[5><2] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[5><2] ) );
  AND2_X1 U448 ( .A1(\warp_gen_fence_regs_wr_cta_id[5><3] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[5><3] ) );
  AND2_X1 U449 ( .A1(\warp_gen_fence_regs_wr_cta_id[6><0] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[6><0] ) );
  AND2_X1 U450 ( .A1(\warp_gen_fence_regs_wr_cta_id[6><1] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[6><1] ) );
  AND2_X1 U451 ( .A1(\warp_gen_fence_regs_wr_cta_id[6><2] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[6><2] ) );
  AND2_X1 U452 ( .A1(\warp_gen_fence_regs_wr_cta_id[6><3] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[6><3] ) );
  AND2_X1 U453 ( .A1(\warp_gen_fence_regs_wr_cta_id[7><0] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[7><0] ) );
  AND2_X1 U454 ( .A1(\warp_gen_fence_regs_wr_cta_id[7><1] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[7><1] ) );
  AND2_X1 U455 ( .A1(\warp_gen_fence_regs_wr_cta_id[7><2] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[7><2] ) );
  AND2_X1 U456 ( .A1(\warp_gen_fence_regs_wr_cta_id[7><3] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[7><3] ) );
  AND2_X1 U457 ( .A1(\warp_gen_fence_regs_wr_cta_id[8><0] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[8><0] ) );
  AND2_X1 U458 ( .A1(\warp_gen_fence_regs_wr_cta_id[8><1] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[8><1] ) );
  AND2_X1 U459 ( .A1(\warp_gen_fence_regs_wr_cta_id[8><2] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[8><2] ) );
  AND2_X1 U460 ( .A1(\warp_gen_fence_regs_wr_cta_id[8><3] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[8><3] ) );
  AND2_X1 U461 ( .A1(\warp_gen_fence_regs_wr_cta_id[9><0] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[9><0] ) );
  AND2_X1 U462 ( .A1(\warp_gen_fence_regs_wr_cta_id[9><1] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[9><1] ) );
  AND2_X1 U463 ( .A1(\warp_gen_fence_regs_wr_cta_id[9><2] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[9><2] ) );
  AND2_X1 U464 ( .A1(\warp_gen_fence_regs_wr_cta_id[9><3] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[9><3] ) );
  AND2_X1 U465 ( .A1(\warp_gen_fence_regs_wr_cta_id[30><0] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[30><0] ) );
  AND2_X1 U466 ( .A1(\warp_gen_fence_regs_wr_cta_id[30><1] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[30><1] ) );
  AND2_X1 U467 ( .A1(\warp_gen_fence_regs_wr_cta_id[30><2] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[30><2] ) );
  AND2_X1 U468 ( .A1(\warp_gen_fence_regs_wr_cta_id[30><3] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[30><3] ) );
  AND2_X1 U469 ( .A1(\warp_gen_fence_regs_wr_cta_id[31><0] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[31><0] ) );
  AND2_X1 U470 ( .A1(\warp_gen_fence_regs_wr_cta_id[31><1] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[31><1] ) );
  AND2_X1 U471 ( .A1(\warp_gen_fence_regs_wr_cta_id[31><2] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[31><2] ) );
  AND2_X1 U472 ( .A1(\warp_gen_fence_regs_wr_cta_id[31><3] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[31><3] ) );
  INV_X1 U473 ( .A(n402), .ZN(n2) );
  INV_X1 U474 ( .A(n391), .ZN(n3) );
  INV_X1 U475 ( .A(n388), .ZN(n4) );
  INV_X1 U476 ( .A(n386), .ZN(n6) );
  INV_X1 U477 ( .A(n385), .ZN(n7) );
  INV_X1 U478 ( .A(n383), .ZN(n9) );
  INV_X1 U479 ( .A(n406), .ZN(n17) );
  INV_X1 U480 ( .A(n405), .ZN(n18) );
  INV_X1 U481 ( .A(n404), .ZN(n19) );
  INV_X1 U482 ( .A(n403), .ZN(n20) );
  INV_X1 U483 ( .A(n400), .ZN(n22) );
  INV_X1 U484 ( .A(n399), .ZN(n23) );
  INV_X1 U485 ( .A(n398), .ZN(n24) );
  INV_X1 U486 ( .A(n397), .ZN(n25) );
  INV_X1 U487 ( .A(n396), .ZN(n26) );
  INV_X1 U488 ( .A(n395), .ZN(n27) );
  INV_X1 U489 ( .A(n392), .ZN(n30) );
  INV_X1 U490 ( .A(n389), .ZN(n32) );
  INV_X1 U491 ( .A(n412), .ZN(n11) );
  INV_X1 U492 ( .A(n410), .ZN(n13) );
  INV_X1 U493 ( .A(n409), .ZN(n14) );
  INV_X1 U494 ( .A(n407), .ZN(n16) );
  INV_X1 U495 ( .A(n413), .ZN(n1) );
  BUF_X1 U496 ( .A(host_reset), .Z(n248) );
  BUF_X1 U497 ( .A(host_reset), .Z(n249) );
  AND2_X1 U498 ( .A1(warp_gen_pool_wr_data[101]), .A2(n176), .ZN(n65) );
  AND2_X1 U499 ( .A1(warp_gen_pool_wr_data[102]), .A2(n176), .ZN(n66) );
  AND2_X1 U500 ( .A1(warp_gen_pool_wr_data[103]), .A2(n176), .ZN(n67) );
  AND2_X1 U501 ( .A1(warp_gen_pool_wr_data[104]), .A2(n176), .ZN(n68) );
  AND2_X1 U502 ( .A1(warp_gen_pool_wr_data[105]), .A2(n176), .ZN(n69) );
  AND2_X1 U503 ( .A1(warp_gen_pool_wr_data[106]), .A2(n176), .ZN(n70) );
  AND2_X1 U504 ( .A1(warp_gen_pool_wr_data[107]), .A2(n176), .ZN(n71) );
  AND2_X1 U505 ( .A1(warp_gen_pool_wr_data[108]), .A2(n176), .ZN(n72) );
  AND2_X1 U506 ( .A1(warp_gen_pool_wr_data[109]), .A2(n176), .ZN(n73) );
  AND2_X1 U507 ( .A1(warp_gen_pool_wr_data[110]), .A2(n176), .ZN(n74) );
  AND2_X1 U508 ( .A1(warp_gen_pool_wr_data[111]), .A2(n176), .ZN(n75) );
  AND2_X1 U509 ( .A1(warp_gen_pool_wr_data[112]), .A2(n176), .ZN(n76) );
  AND2_X1 U510 ( .A1(warp_gen_pool_wr_data[113]), .A2(n176), .ZN(n77) );
  AND2_X1 U511 ( .A1(warp_gen_pool_wr_data[114]), .A2(n176), .ZN(n78) );
  AND2_X1 U512 ( .A1(warp_gen_pool_wr_data[115]), .A2(n176), .ZN(n79) );
  AND2_X1 U513 ( .A1(warp_gen_pool_wr_data[116]), .A2(n176), .ZN(n80) );
  INV_X1 U514 ( .A(n208), .ZN(n251) );
  AOI22_X1 U515 ( .A1(n164), .A2(warp_gen_state_wr_en), .B1(
        warp_sched_state_wr_en), .B2(n181), .ZN(n208) );
  INV_X1 U516 ( .A(n214), .ZN(n260) );
  AOI22_X1 U517 ( .A1(warp_gen_state_addr[1]), .A2(n163), .B1(
        warp_sched_state_addr[1]), .B2(n179), .ZN(n214) );
  INV_X1 U518 ( .A(n213), .ZN(n254) );
  AOI22_X1 U519 ( .A1(warp_gen_state_addr[2]), .A2(n163), .B1(
        warp_sched_state_addr[2]), .B2(n179), .ZN(n213) );
  INV_X1 U520 ( .A(n346), .ZN(n253) );
  AOI22_X1 U521 ( .A1(warp_gen_pool_addr[3]), .A2(n163), .B1(
        warp_sched_pool_addr[3]), .B2(n180), .ZN(n346) );
  INV_X1 U522 ( .A(n345), .ZN(n259) );
  AOI22_X1 U523 ( .A1(warp_gen_pool_addr[4]), .A2(n163), .B1(
        warp_sched_pool_addr[4]), .B2(n180), .ZN(n345) );
  INV_X1 U524 ( .A(n215), .ZN(n256) );
  AOI22_X1 U525 ( .A1(warp_gen_state_addr[0]), .A2(n164), .B1(
        warp_sched_state_addr[0]), .B2(n180), .ZN(n215) );
  INV_X1 U526 ( .A(n212), .ZN(n252) );
  AOI22_X1 U527 ( .A1(warp_gen_state_addr[3]), .A2(n164), .B1(
        warp_sched_state_addr[3]), .B2(n179), .ZN(n212) );
  INV_X1 U528 ( .A(n211), .ZN(n258) );
  AOI22_X1 U529 ( .A1(warp_gen_state_addr[4]), .A2(n164), .B1(
        warp_sched_state_addr[4]), .B2(n179), .ZN(n211) );
  INV_X1 U530 ( .A(n349), .ZN(n257) );
  AOI22_X1 U531 ( .A1(warp_gen_pool_addr[0]), .A2(n164), .B1(
        warp_sched_pool_addr[0]), .B2(n181), .ZN(n349) );
  INV_X1 U532 ( .A(n348), .ZN(n261) );
  AOI22_X1 U533 ( .A1(warp_gen_pool_addr[1]), .A2(n164), .B1(
        warp_sched_pool_addr[1]), .B2(n181), .ZN(n348) );
  INV_X1 U534 ( .A(n347), .ZN(n255) );
  AOI22_X1 U535 ( .A1(warp_gen_pool_addr[2]), .A2(n164), .B1(
        warp_sched_pool_addr[2]), .B2(n180), .ZN(n347) );
  AND2_X1 U536 ( .A1(warp_gen_pool_wr_data[0]), .A2(n175), .ZN(n81) );
  AND2_X1 U537 ( .A1(warp_gen_pool_wr_data[117]), .A2(n175), .ZN(n82) );
  AND2_X1 U538 ( .A1(warp_gen_pool_wr_data[118]), .A2(n175), .ZN(n83) );
  AND2_X1 U539 ( .A1(warp_gen_pool_wr_data[119]), .A2(n175), .ZN(n84) );
  AND2_X1 U540 ( .A1(warp_gen_pool_wr_data[120]), .A2(n175), .ZN(n85) );
  AND2_X1 U541 ( .A1(warp_gen_pool_wr_data[121]), .A2(n175), .ZN(n86) );
  AND2_X1 U542 ( .A1(warp_gen_pool_wr_data[122]), .A2(n175), .ZN(n87) );
  AND2_X1 U543 ( .A1(warp_gen_pool_wr_data[123]), .A2(n175), .ZN(n88) );
  AND2_X1 U544 ( .A1(warp_gen_pool_wr_en), .A2(n178), .ZN(n89) );
  AND2_X1 U545 ( .A1(warp_gen_pool_wr_data[37]), .A2(n177), .ZN(n90) );
  AND2_X1 U546 ( .A1(warp_gen_pool_wr_data[38]), .A2(n178), .ZN(n91) );
  AND2_X1 U547 ( .A1(warp_gen_pool_wr_data[39]), .A2(n176), .ZN(n92) );
  AND2_X1 U548 ( .A1(warp_gen_pool_wr_data[40]), .A2(n178), .ZN(n93) );
  AND2_X1 U549 ( .A1(warp_gen_pool_wr_data[41]), .A2(n177), .ZN(n94) );
  AND2_X1 U550 ( .A1(warp_gen_pool_wr_data[42]), .A2(n177), .ZN(n95) );
  AND2_X1 U551 ( .A1(warp_gen_pool_wr_data[43]), .A2(n176), .ZN(n96) );
  AND2_X1 U552 ( .A1(warp_gen_pool_wr_data[44]), .A2(n178), .ZN(n97) );
  AND2_X1 U553 ( .A1(warp_gen_pool_wr_data[45]), .A2(n177), .ZN(n98) );
  AND2_X1 U554 ( .A1(warp_gen_pool_wr_data[46]), .A2(n176), .ZN(n99) );
  AND2_X1 U555 ( .A1(warp_gen_pool_wr_data[47]), .A2(n176), .ZN(n100) );
  AND2_X1 U556 ( .A1(warp_gen_pool_wr_data[48]), .A2(n178), .ZN(n101) );
  AND2_X1 U557 ( .A1(warp_gen_pool_wr_data[49]), .A2(n177), .ZN(n102) );
  AND2_X1 U558 ( .A1(warp_gen_pool_wr_data[50]), .A2(n178), .ZN(n103) );
  AND2_X1 U559 ( .A1(warp_gen_pool_wr_data[51]), .A2(n176), .ZN(n104) );
  AND2_X1 U560 ( .A1(warp_gen_pool_wr_data[5]), .A2(n178), .ZN(n105) );
  AND2_X1 U561 ( .A1(warp_gen_pool_wr_data[6]), .A2(n178), .ZN(n106) );
  AND2_X1 U562 ( .A1(warp_gen_pool_wr_data[7]), .A2(n178), .ZN(n107) );
  AND2_X1 U563 ( .A1(warp_gen_pool_wr_data[8]), .A2(n178), .ZN(n108) );
  AND2_X1 U564 ( .A1(warp_gen_pool_wr_data[9]), .A2(n178), .ZN(n109) );
  AND2_X1 U565 ( .A1(warp_gen_pool_wr_data[10]), .A2(n178), .ZN(n110) );
  AND2_X1 U566 ( .A1(warp_gen_pool_wr_data[11]), .A2(n178), .ZN(n111) );
  AND2_X1 U567 ( .A1(warp_gen_pool_wr_data[12]), .A2(n178), .ZN(n112) );
  AND2_X1 U568 ( .A1(warp_gen_pool_wr_data[13]), .A2(n178), .ZN(n113) );
  AND2_X1 U569 ( .A1(warp_gen_pool_wr_data[14]), .A2(n178), .ZN(n114) );
  AND2_X1 U570 ( .A1(warp_gen_pool_wr_data[15]), .A2(n178), .ZN(n115) );
  AND2_X1 U571 ( .A1(warp_gen_pool_wr_data[16]), .A2(n178), .ZN(n116) );
  AND2_X1 U572 ( .A1(warp_gen_pool_wr_data[17]), .A2(n178), .ZN(n117) );
  AND2_X1 U573 ( .A1(warp_gen_pool_wr_data[18]), .A2(n178), .ZN(n118) );
  AND2_X1 U574 ( .A1(warp_gen_pool_wr_data[19]), .A2(n178), .ZN(n119) );
  AND2_X1 U575 ( .A1(warp_gen_pool_wr_data[20]), .A2(n178), .ZN(n120) );
  AND2_X1 U576 ( .A1(warp_gen_pool_wr_data[21]), .A2(n177), .ZN(n121) );
  AND2_X1 U577 ( .A1(warp_gen_pool_wr_data[22]), .A2(n177), .ZN(n122) );
  AND2_X1 U578 ( .A1(warp_gen_pool_wr_data[23]), .A2(n177), .ZN(n123) );
  AND2_X1 U579 ( .A1(warp_gen_pool_wr_data[24]), .A2(n177), .ZN(n124) );
  AND2_X1 U580 ( .A1(warp_gen_pool_wr_data[25]), .A2(n177), .ZN(n125) );
  AND2_X1 U581 ( .A1(warp_gen_pool_wr_data[26]), .A2(n177), .ZN(n126) );
  AND2_X1 U582 ( .A1(warp_gen_pool_wr_data[27]), .A2(n177), .ZN(n127) );
  AND2_X1 U583 ( .A1(warp_gen_pool_wr_data[28]), .A2(n177), .ZN(n128) );
  AND2_X1 U584 ( .A1(warp_gen_pool_wr_data[29]), .A2(n177), .ZN(n129) );
  AND2_X1 U585 ( .A1(warp_gen_pool_wr_data[30]), .A2(n177), .ZN(n130) );
  AND2_X1 U586 ( .A1(warp_gen_pool_wr_data[31]), .A2(n177), .ZN(n131) );
  AND2_X1 U587 ( .A1(warp_gen_pool_wr_data[32]), .A2(n177), .ZN(n132) );
  AND2_X1 U588 ( .A1(warp_gen_pool_wr_data[33]), .A2(n177), .ZN(n133) );
  AND2_X1 U589 ( .A1(warp_gen_pool_wr_data[34]), .A2(n177), .ZN(n134) );
  AND2_X1 U590 ( .A1(warp_gen_pool_wr_data[35]), .A2(n177), .ZN(n135) );
  AND2_X1 U591 ( .A1(warp_gen_pool_wr_data[36]), .A2(n177), .ZN(n136) );
  AND2_X1 U592 ( .A1(warp_gen_pool_wr_data[52]), .A2(n176), .ZN(n137) );
  AND2_X1 U593 ( .A1(warp_gen_pool_wr_data[53]), .A2(n178), .ZN(n138) );
  AND2_X1 U594 ( .A1(warp_gen_pool_wr_data[54]), .A2(n177), .ZN(n139) );
  AND2_X1 U595 ( .A1(warp_gen_pool_wr_data[55]), .A2(n176), .ZN(n140) );
  AND2_X1 U596 ( .A1(warp_gen_pool_wr_data[56]), .A2(n178), .ZN(n141) );
  AND2_X1 U597 ( .A1(warp_gen_pool_wr_data[57]), .A2(n177), .ZN(n142) );
  AND2_X1 U598 ( .A1(warp_gen_pool_wr_data[58]), .A2(n176), .ZN(n143) );
  AND2_X1 U599 ( .A1(warp_gen_pool_wr_data[59]), .A2(n178), .ZN(n144) );
  AND2_X1 U600 ( .A1(warp_gen_pool_wr_data[60]), .A2(n177), .ZN(n145) );
  AND2_X1 U601 ( .A1(warp_gen_pool_wr_data[61]), .A2(n176), .ZN(n146) );
  AND2_X1 U602 ( .A1(warp_gen_pool_wr_data[62]), .A2(n178), .ZN(n147) );
  AND2_X1 U603 ( .A1(warp_gen_pool_wr_data[63]), .A2(n177), .ZN(n148) );
  AND2_X1 U604 ( .A1(warp_gen_pool_wr_data[97]), .A2(n176), .ZN(n149) );
  AND2_X1 U605 ( .A1(warp_gen_pool_wr_data[98]), .A2(n178), .ZN(n150) );
  AND2_X1 U606 ( .A1(warp_gen_pool_wr_data[99]), .A2(n177), .ZN(n151) );
  AND2_X1 U607 ( .A1(warp_gen_pool_wr_data[100]), .A2(n176), .ZN(n152) );
  AND2_X1 U608 ( .A1(warp_gen_pool_wr_data[1]), .A2(n178), .ZN(n153) );
  AND2_X1 U609 ( .A1(warp_gen_pool_wr_data[2]), .A2(n177), .ZN(n154) );
  AND2_X1 U610 ( .A1(warp_gen_pool_wr_data[3]), .A2(n177), .ZN(n155) );
  AND2_X1 U611 ( .A1(warp_gen_pool_wr_data[4]), .A2(n176), .ZN(n156) );
  AND2_X1 U612 ( .A1(\warp_sched_state_wr_data[0] ), .A2(n224), .ZN(n157) );
  INV_X1 U613 ( .A(n220), .ZN(n161) );
  INV_X1 U614 ( .A(n220), .ZN(n162) );
  INV_X1 U615 ( .A(n219), .ZN(n166) );
  INV_X1 U616 ( .A(n220), .ZN(n168) );
  INV_X1 U617 ( .A(n219), .ZN(n169) );
  INV_X1 U618 ( .A(n221), .ZN(n173) );
  INV_X1 U619 ( .A(n221), .ZN(n176) );
endmodule




module warps_done_lut ( clk_in, host_reset, num_warps_in, warps_done_mask );
  input [4:0] num_warps_in;
  output [31:0] warps_done_mask;
  input clk_in, host_reset;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n69, n70, n71;

  DFFR_X1 \warps_done_mask_reg[31]  ( .D(n68), .CK(clk_in), .RN(n10), .Q(
        warps_done_mask[31]) );
  DFFR_X1 \warps_done_mask_reg[30]  ( .D(n67), .CK(clk_in), .RN(n9), .Q(
        warps_done_mask[30]) );
  DFFR_X1 \warps_done_mask_reg[29]  ( .D(n21), .CK(clk_in), .RN(n9), .Q(
        warps_done_mask[29]) );
  DFFR_X1 \warps_done_mask_reg[28]  ( .D(n66), .CK(clk_in), .RN(n9), .Q(
        warps_done_mask[28]) );
  DFFR_X1 \warps_done_mask_reg[27]  ( .D(n22), .CK(clk_in), .RN(n9), .Q(
        warps_done_mask[27]) );
  DFFR_X1 \warps_done_mask_reg[26]  ( .D(n65), .CK(clk_in), .RN(n9), .Q(
        warps_done_mask[26]) );
  DFFR_X1 \warps_done_mask_reg[25]  ( .D(n23), .CK(clk_in), .RN(n9), .Q(
        warps_done_mask[25]) );
  DFFR_X1 \warps_done_mask_reg[24]  ( .D(n64), .CK(clk_in), .RN(n9), .Q(
        warps_done_mask[24]) );
  DFFR_X1 \warps_done_mask_reg[23]  ( .D(n24), .CK(clk_in), .RN(n9), .Q(
        warps_done_mask[23]) );
  DFFR_X1 \warps_done_mask_reg[22]  ( .D(n63), .CK(clk_in), .RN(n9), .Q(
        warps_done_mask[22]) );
  DFFR_X1 \warps_done_mask_reg[21]  ( .D(n25), .CK(clk_in), .RN(n9), .Q(
        warps_done_mask[21]) );
  DFFR_X1 \warps_done_mask_reg[20]  ( .D(n62), .CK(clk_in), .RN(n9), .Q(
        warps_done_mask[20]) );
  DFFR_X1 \warps_done_mask_reg[19]  ( .D(n26), .CK(clk_in), .RN(n10), .Q(
        warps_done_mask[19]) );
  DFFR_X1 \warps_done_mask_reg[18]  ( .D(n61), .CK(clk_in), .RN(n10), .Q(
        warps_done_mask[18]) );
  DFFR_X1 \warps_done_mask_reg[17]  ( .D(n13), .CK(clk_in), .RN(n10), .Q(
        warps_done_mask[17]) );
  DFFR_X1 \warps_done_mask_reg[16]  ( .D(n60), .CK(clk_in), .RN(n10), .Q(
        warps_done_mask[16]) );
  SDFFR_X1 \warps_done_mask_reg[15]  ( .D(n13), .SI(1'b1), .SE(num_warps_in[4]), .CK(clk_in), .RN(n11), .Q(warps_done_mask[15]) );
  DFFR_X1 \warps_done_mask_reg[14]  ( .D(n14), .CK(clk_in), .RN(n10), .Q(
        warps_done_mask[14]) );
  SDFFR_X1 \warps_done_mask_reg[13]  ( .D(n59), .SI(1'b1), .SE(n43), .CK(
        clk_in), .RN(n11), .Q(warps_done_mask[13]) );
  DFFR_X1 \warps_done_mask_reg[12]  ( .D(n15), .CK(clk_in), .RN(n10), .Q(
        warps_done_mask[12]) );
  SDFFR_X1 \warps_done_mask_reg[11]  ( .D(n58), .SI(1'b1), .SE(n70), .CK(
        clk_in), .RN(n11), .Q(warps_done_mask[11]) );
  DFFR_X1 \warps_done_mask_reg[10]  ( .D(n16), .CK(clk_in), .RN(n10), .Q(
        warps_done_mask[10]) );
  SDFFR_X1 \warps_done_mask_reg[9]  ( .D(n57), .SI(1'b1), .SE(n31), .CK(clk_in), .RN(n11), .Q(warps_done_mask[9]) );
  DFFR_X1 \warps_done_mask_reg[8]  ( .D(n17), .CK(clk_in), .RN(n10), .Q(
        warps_done_mask[8]) );
  SDFFR_X1 \warps_done_mask_reg[7]  ( .D(n56), .SI(1'b1), .SE(num_warps_in[3]), 
        .CK(clk_in), .RN(n11), .Q(warps_done_mask[7]) );
  DFFR_X1 \warps_done_mask_reg[6]  ( .D(n18), .CK(clk_in), .RN(n10), .Q(
        warps_done_mask[6]) );
  SDFFR_X1 \warps_done_mask_reg[5]  ( .D(n55), .SI(1'b1), .SE(n30), .CK(clk_in), .RN(n11), .Q(warps_done_mask[5]) );
  DFFR_X1 \warps_done_mask_reg[4]  ( .D(n19), .CK(clk_in), .RN(n10), .Q(
        warps_done_mask[4]) );
  SDFFR_X1 \warps_done_mask_reg[3]  ( .D(n54), .SI(1'b1), .SE(num_warps_in[2]), 
        .CK(clk_in), .RN(n11), .Q(warps_done_mask[3]) );
  DFFR_X1 \warps_done_mask_reg[2]  ( .D(n20), .CK(clk_in), .RN(n10), .Q(
        warps_done_mask[2]) );
  SDFFR_X1 \warps_done_mask_reg[1]  ( .D(n53), .SI(1'b1), .SE(num_warps_in[1]), 
        .CK(clk_in), .RN(n11), .Q(warps_done_mask[1]) );
  DFFR_X1 \warps_done_mask_reg[0]  ( .D(1'b1), .CK(clk_in), .RN(n9), .Q(
        warps_done_mask[0]) );
  NAND2_X1 U60 ( .A1(n34), .A2(n69), .ZN(n53) );
  NAND2_X1 U61 ( .A1(n35), .A2(n36), .ZN(n54) );
  NAND2_X1 U62 ( .A1(n37), .A2(n71), .ZN(n55) );
  NAND2_X1 U63 ( .A1(n38), .A2(n39), .ZN(n56) );
  NAND2_X1 U64 ( .A1(n40), .A2(n41), .ZN(n57) );
  NAND2_X1 U65 ( .A1(n27), .A2(n42), .ZN(n58) );
  NAND2_X1 U66 ( .A1(n44), .A2(n45), .ZN(n60) );
  NAND2_X1 U67 ( .A1(num_warps_in[2]), .A2(num_warps_in[1]), .ZN(n35) );
  NAND2_X1 U68 ( .A1(num_warps_in[3]), .A2(num_warps_in[1]), .ZN(n38) );
  NAND2_X1 U69 ( .A1(num_warps_in[3]), .A2(num_warps_in[2]), .ZN(n40) );
  NAND2_X1 U70 ( .A1(num_warps_in[4]), .A2(num_warps_in[0]), .ZN(n44) );
  INV_X1 U11 ( .A(n43), .ZN(n27) );
  BUF_X1 U12 ( .A(n12), .Z(n9) );
  BUF_X1 U13 ( .A(n12), .Z(n10) );
  BUF_X1 U14 ( .A(n12), .Z(n11) );
  NOR3_X1 U15 ( .A1(n69), .A2(n28), .A3(n71), .ZN(n43) );
  OAI21_X1 U16 ( .B1(n44), .B2(n35), .A(n48), .ZN(n63) );
  OAI21_X1 U17 ( .B1(n44), .B2(n38), .A(n50), .ZN(n65) );
  OAI21_X1 U18 ( .B1(n44), .B2(n40), .A(n51), .ZN(n66) );
  OAI21_X1 U19 ( .B1(n44), .B2(n27), .A(n29), .ZN(n67) );
  INV_X1 U20 ( .A(n68), .ZN(n29) );
  OAI21_X1 U21 ( .B1(n28), .B2(n44), .A(n46), .ZN(n61) );
  OAI21_X1 U22 ( .B1(n69), .B2(n44), .A(n47), .ZN(n62) );
  OAI21_X1 U23 ( .B1(n71), .B2(n44), .A(n49), .ZN(n64) );
  INV_X1 U24 ( .A(n40), .ZN(n70) );
  INV_X1 U25 ( .A(n36), .ZN(n18) );
  INV_X1 U26 ( .A(n34), .ZN(n19) );
  INV_X1 U27 ( .A(n35), .ZN(n30) );
  INV_X1 U28 ( .A(n38), .ZN(n31) );
  INV_X1 U29 ( .A(n45), .ZN(n13) );
  INV_X1 U30 ( .A(n47), .ZN(n25) );
  INV_X1 U31 ( .A(n39), .ZN(n16) );
  INV_X1 U32 ( .A(n41), .ZN(n15) );
  INV_X1 U33 ( .A(n42), .ZN(n14) );
  INV_X1 U34 ( .A(n46), .ZN(n26) );
  INV_X1 U35 ( .A(n48), .ZN(n24) );
  INV_X1 U36 ( .A(n37), .ZN(n17) );
  INV_X1 U37 ( .A(n49), .ZN(n23) );
  INV_X1 U38 ( .A(n50), .ZN(n22) );
  INV_X1 U39 ( .A(n51), .ZN(n21) );
  INV_X1 U40 ( .A(host_reset), .ZN(n12) );
  AOI21_X1 U41 ( .B1(num_warps_in[2]), .B2(num_warps_in[4]), .A(n62), .ZN(n46)
         );
  AOI21_X1 U42 ( .B1(num_warps_in[3]), .B2(num_warps_in[4]), .A(n64), .ZN(n48)
         );
  AOI21_X1 U43 ( .B1(num_warps_in[4]), .B2(n30), .A(n63), .ZN(n47) );
  AOI21_X1 U44 ( .B1(num_warps_in[4]), .B2(n31), .A(n65), .ZN(n49) );
  AOI21_X1 U45 ( .B1(num_warps_in[4]), .B2(n70), .A(n66), .ZN(n50) );
  AOI21_X1 U46 ( .B1(num_warps_in[4]), .B2(n43), .A(n67), .ZN(n51) );
  AOI21_X1 U47 ( .B1(num_warps_in[1]), .B2(num_warps_in[4]), .A(n61), .ZN(n45)
         );
  AOI21_X1 U48 ( .B1(num_warps_in[2]), .B2(num_warps_in[0]), .A(n54), .ZN(n34)
         );
  AOI21_X1 U49 ( .B1(num_warps_in[3]), .B2(num_warps_in[0]), .A(n56), .ZN(n37)
         );
  AOI21_X1 U50 ( .B1(num_warps_in[0]), .B2(n30), .A(n55), .ZN(n36) );
  AOI21_X1 U51 ( .B1(num_warps_in[0]), .B2(n31), .A(n57), .ZN(n39) );
  AOI21_X1 U52 ( .B1(num_warps_in[0]), .B2(n70), .A(n58), .ZN(n41) );
  AOI21_X1 U53 ( .B1(num_warps_in[0]), .B2(n43), .A(n59), .ZN(n42) );
  INV_X1 U54 ( .A(num_warps_in[3]), .ZN(n71) );
  INV_X1 U55 ( .A(num_warps_in[2]), .ZN(n69) );
  INV_X1 U56 ( .A(num_warps_in[1]), .ZN(n28) );
  OR2_X1 U57 ( .A1(n60), .A2(num_warps_in[4]), .ZN(n59) );
  NOR4_X1 U58 ( .A1(num_warps_in[0]), .A2(num_warps_in[1]), .A3(n52), .A4(
        num_warps_in[2]), .ZN(n68) );
  OR2_X1 U71 ( .A1(num_warps_in[4]), .A2(num_warps_in[3]), .ZN(n52) );
  INV_X1 U72 ( .A(n33), .ZN(n20) );
  AOI21_X1 U73 ( .B1(num_warps_in[1]), .B2(num_warps_in[0]), .A(n53), .ZN(n33)
         );
endmodule












