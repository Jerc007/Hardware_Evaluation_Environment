

module warp_unit ( clk_in, host_reset, warp_scheduler_reset, 
        warp_generator_en, pipeline_write_done, pipeline_stall_in, 
        threads_per_block_in, num_blocks_in, warps_per_block_in, 
        shared_mem_base_addr_in, shared_mem_size_in, gprs_size_in, block_x_in, 
        block_y_in, block_z_in, grid_x_in, grid_y_in, block_idx_in, warp_id_in, 
        warp_lane_id_in, cta_id_in, initial_mask_in, current_mask_in, 
        shmem_base_addr_in, gprs_base_addr_in, next_pc_in, warp_state_in, 
        program_cntr_out, warp_id_out, warp_lane_id_out, cta_id_out, 
        initial_mask_out, current_mask_out, shmem_base_addr_out, gprs_size_out, 
        gprs_base_addr_out, num_warps_out, warp_generator_done, 
        pipeline_stall_out, warp_scheduler_done, pipeline_warpunit_done, 
        fetch_en );
  input [11:0] threads_per_block_in;
  input [3:0] num_blocks_in;
  input [5:0] warps_per_block_in;
  input [31:0] shared_mem_base_addr_in;
  input [31:0] shared_mem_size_in;
  input [8:0] gprs_size_in;
  input [15:0] block_x_in;
  input [15:0] block_y_in;
  input [15:0] block_z_in;
  input [15:0] grid_x_in;
  input [15:0] grid_y_in;
  input [15:0] block_idx_in;
  input [4:0] warp_id_in;
  input [1:0] warp_lane_id_in;
  input [3:0] cta_id_in;
  input [31:0] initial_mask_in;
  input [31:0] current_mask_in;
  input [13:0] shmem_base_addr_in;
  input [8:0] gprs_base_addr_in;
  input [31:0] next_pc_in;
  input [1:0] warp_state_in;
  output [31:0] program_cntr_out;
  output [4:0] warp_id_out;
  output [1:0] warp_lane_id_out;
  output [3:0] cta_id_out;
  output [31:0] initial_mask_out;
  output [31:0] current_mask_out;
  output [13:0] shmem_base_addr_out;
  output [8:0] gprs_size_out;
  output [8:0] gprs_base_addr_out;
  output [4:0] num_warps_out;
  input clk_in, host_reset, warp_scheduler_reset, warp_generator_en,
         pipeline_write_done, pipeline_stall_in;
  output warp_generator_done, pipeline_stall_out, warp_scheduler_done,
         pipeline_warpunit_done, fetch_en;
  wire   warp_gen_pool_wr_en, warp_gen_state_wr_en,
         \warp_gen_fence_regs_wr_cta_id[31><3] ,
         \warp_gen_fence_regs_wr_cta_id[31><2] ,
         \warp_gen_fence_regs_wr_cta_id[31><1] ,
         \warp_gen_fence_regs_wr_cta_id[31><0] ,
         \warp_gen_fence_regs_wr_cta_id[30><3] ,
         \warp_gen_fence_regs_wr_cta_id[30><2] ,
         \warp_gen_fence_regs_wr_cta_id[30><1] ,
         \warp_gen_fence_regs_wr_cta_id[30><0] ,
         \warp_gen_fence_regs_wr_cta_id[29><3] ,
         \warp_gen_fence_regs_wr_cta_id[29><2] ,
         \warp_gen_fence_regs_wr_cta_id[29><1] ,
         \warp_gen_fence_regs_wr_cta_id[29><0] ,
         \warp_gen_fence_regs_wr_cta_id[28><3] ,
         \warp_gen_fence_regs_wr_cta_id[28><2] ,
         \warp_gen_fence_regs_wr_cta_id[28><1] ,
         \warp_gen_fence_regs_wr_cta_id[28><0] ,
         \warp_gen_fence_regs_wr_cta_id[27><3] ,
         \warp_gen_fence_regs_wr_cta_id[27><2] ,
         \warp_gen_fence_regs_wr_cta_id[27><1] ,
         \warp_gen_fence_regs_wr_cta_id[27><0] ,
         \warp_gen_fence_regs_wr_cta_id[26><3] ,
         \warp_gen_fence_regs_wr_cta_id[26><2] ,
         \warp_gen_fence_regs_wr_cta_id[26><1] ,
         \warp_gen_fence_regs_wr_cta_id[26><0] ,
         \warp_gen_fence_regs_wr_cta_id[25><3] ,
         \warp_gen_fence_regs_wr_cta_id[25><2] ,
         \warp_gen_fence_regs_wr_cta_id[25><1] ,
         \warp_gen_fence_regs_wr_cta_id[25><0] ,
         \warp_gen_fence_regs_wr_cta_id[24><3] ,
         \warp_gen_fence_regs_wr_cta_id[24><2] ,
         \warp_gen_fence_regs_wr_cta_id[24><1] ,
         \warp_gen_fence_regs_wr_cta_id[24><0] ,
         \warp_gen_fence_regs_wr_cta_id[23><3] ,
         \warp_gen_fence_regs_wr_cta_id[23><2] ,
         \warp_gen_fence_regs_wr_cta_id[23><1] ,
         \warp_gen_fence_regs_wr_cta_id[23><0] ,
         \warp_gen_fence_regs_wr_cta_id[22><3] ,
         \warp_gen_fence_regs_wr_cta_id[22><2] ,
         \warp_gen_fence_regs_wr_cta_id[22><1] ,
         \warp_gen_fence_regs_wr_cta_id[22><0] ,
         \warp_gen_fence_regs_wr_cta_id[21><3] ,
         \warp_gen_fence_regs_wr_cta_id[21><2] ,
         \warp_gen_fence_regs_wr_cta_id[21><1] ,
         \warp_gen_fence_regs_wr_cta_id[21><0] ,
         \warp_gen_fence_regs_wr_cta_id[20><3] ,
         \warp_gen_fence_regs_wr_cta_id[20><2] ,
         \warp_gen_fence_regs_wr_cta_id[20><1] ,
         \warp_gen_fence_regs_wr_cta_id[20><0] ,
         \warp_gen_fence_regs_wr_cta_id[19><3] ,
         \warp_gen_fence_regs_wr_cta_id[19><2] ,
         \warp_gen_fence_regs_wr_cta_id[19><1] ,
         \warp_gen_fence_regs_wr_cta_id[19><0] ,
         \warp_gen_fence_regs_wr_cta_id[18><3] ,
         \warp_gen_fence_regs_wr_cta_id[18><2] ,
         \warp_gen_fence_regs_wr_cta_id[18><1] ,
         \warp_gen_fence_regs_wr_cta_id[18><0] ,
         \warp_gen_fence_regs_wr_cta_id[17><3] ,
         \warp_gen_fence_regs_wr_cta_id[17><2] ,
         \warp_gen_fence_regs_wr_cta_id[17><1] ,
         \warp_gen_fence_regs_wr_cta_id[17><0] ,
         \warp_gen_fence_regs_wr_cta_id[16><3] ,
         \warp_gen_fence_regs_wr_cta_id[16><2] ,
         \warp_gen_fence_regs_wr_cta_id[16><1] ,
         \warp_gen_fence_regs_wr_cta_id[16><0] ,
         \warp_gen_fence_regs_wr_cta_id[15><3] ,
         \warp_gen_fence_regs_wr_cta_id[15><2] ,
         \warp_gen_fence_regs_wr_cta_id[15><1] ,
         \warp_gen_fence_regs_wr_cta_id[15><0] ,
         \warp_gen_fence_regs_wr_cta_id[14><3] ,
         \warp_gen_fence_regs_wr_cta_id[14><2] ,
         \warp_gen_fence_regs_wr_cta_id[14><1] ,
         \warp_gen_fence_regs_wr_cta_id[14><0] ,
         \warp_gen_fence_regs_wr_cta_id[13><3] ,
         \warp_gen_fence_regs_wr_cta_id[13><2] ,
         \warp_gen_fence_regs_wr_cta_id[13><1] ,
         \warp_gen_fence_regs_wr_cta_id[13><0] ,
         \warp_gen_fence_regs_wr_cta_id[12><3] ,
         \warp_gen_fence_regs_wr_cta_id[12><2] ,
         \warp_gen_fence_regs_wr_cta_id[12><1] ,
         \warp_gen_fence_regs_wr_cta_id[12><0] ,
         \warp_gen_fence_regs_wr_cta_id[11><3] ,
         \warp_gen_fence_regs_wr_cta_id[11><2] ,
         \warp_gen_fence_regs_wr_cta_id[11><1] ,
         \warp_gen_fence_regs_wr_cta_id[11><0] ,
         \warp_gen_fence_regs_wr_cta_id[10><3] ,
         \warp_gen_fence_regs_wr_cta_id[10><2] ,
         \warp_gen_fence_regs_wr_cta_id[10><1] ,
         \warp_gen_fence_regs_wr_cta_id[10><0] ,
         \warp_gen_fence_regs_wr_cta_id[9><3] ,
         \warp_gen_fence_regs_wr_cta_id[9><2] ,
         \warp_gen_fence_regs_wr_cta_id[9><1] ,
         \warp_gen_fence_regs_wr_cta_id[9><0] ,
         \warp_gen_fence_regs_wr_cta_id[8><3] ,
         \warp_gen_fence_regs_wr_cta_id[8><2] ,
         \warp_gen_fence_regs_wr_cta_id[8><1] ,
         \warp_gen_fence_regs_wr_cta_id[8><0] ,
         \warp_gen_fence_regs_wr_cta_id[7><3] ,
         \warp_gen_fence_regs_wr_cta_id[7><2] ,
         \warp_gen_fence_regs_wr_cta_id[7><1] ,
         \warp_gen_fence_regs_wr_cta_id[7><0] ,
         \warp_gen_fence_regs_wr_cta_id[6><3] ,
         \warp_gen_fence_regs_wr_cta_id[6><2] ,
         \warp_gen_fence_regs_wr_cta_id[6><1] ,
         \warp_gen_fence_regs_wr_cta_id[6><0] ,
         \warp_gen_fence_regs_wr_cta_id[5><3] ,
         \warp_gen_fence_regs_wr_cta_id[5><2] ,
         \warp_gen_fence_regs_wr_cta_id[5><1] ,
         \warp_gen_fence_regs_wr_cta_id[5><0] ,
         \warp_gen_fence_regs_wr_cta_id[4><3] ,
         \warp_gen_fence_regs_wr_cta_id[4><2] ,
         \warp_gen_fence_regs_wr_cta_id[4><1] ,
         \warp_gen_fence_regs_wr_cta_id[4><0] ,
         \warp_gen_fence_regs_wr_cta_id[3><3] ,
         \warp_gen_fence_regs_wr_cta_id[3><2] ,
         \warp_gen_fence_regs_wr_cta_id[3><1] ,
         \warp_gen_fence_regs_wr_cta_id[3><0] ,
         \warp_gen_fence_regs_wr_cta_id[2><3] ,
         \warp_gen_fence_regs_wr_cta_id[2><2] ,
         \warp_gen_fence_regs_wr_cta_id[2><1] ,
         \warp_gen_fence_regs_wr_cta_id[2><0] ,
         \warp_gen_fence_regs_wr_cta_id[1><3] ,
         \warp_gen_fence_regs_wr_cta_id[1><2] ,
         \warp_gen_fence_regs_wr_cta_id[1><1] ,
         \warp_gen_fence_regs_wr_cta_id[1><0] ,
         \warp_gen_fence_regs_wr_cta_id[0><3] ,
         \warp_gen_fence_regs_wr_cta_id[0><2] ,
         \warp_gen_fence_regs_wr_cta_id[0><1] ,
         \warp_gen_fence_regs_wr_cta_id[0><0] , warp_sched_state_wr_en,
         \warp_sched_state_wr_data[0] , warp_pool_wr_en_b, warp_state_wr_en_b,
         \warp_checker_fence_regs_rd_cta_id[31><3] ,
         \warp_checker_fence_regs_rd_cta_id[31><2] ,
         \warp_checker_fence_regs_rd_cta_id[31><1] ,
         \warp_checker_fence_regs_rd_cta_id[31><0] ,
         \warp_checker_fence_regs_rd_cta_id[30><3] ,
         \warp_checker_fence_regs_rd_cta_id[30><2] ,
         \warp_checker_fence_regs_rd_cta_id[30><1] ,
         \warp_checker_fence_regs_rd_cta_id[30><0] ,
         \warp_checker_fence_regs_rd_cta_id[29><3] ,
         \warp_checker_fence_regs_rd_cta_id[29><2] ,
         \warp_checker_fence_regs_rd_cta_id[29><1] ,
         \warp_checker_fence_regs_rd_cta_id[29><0] ,
         \warp_checker_fence_regs_rd_cta_id[28><3] ,
         \warp_checker_fence_regs_rd_cta_id[28><2] ,
         \warp_checker_fence_regs_rd_cta_id[28><1] ,
         \warp_checker_fence_regs_rd_cta_id[28><0] ,
         \warp_checker_fence_regs_rd_cta_id[27><3] ,
         \warp_checker_fence_regs_rd_cta_id[27><2] ,
         \warp_checker_fence_regs_rd_cta_id[27><1] ,
         \warp_checker_fence_regs_rd_cta_id[27><0] ,
         \warp_checker_fence_regs_rd_cta_id[26><3] ,
         \warp_checker_fence_regs_rd_cta_id[26><2] ,
         \warp_checker_fence_regs_rd_cta_id[26><1] ,
         \warp_checker_fence_regs_rd_cta_id[26><0] ,
         \warp_checker_fence_regs_rd_cta_id[25><3] ,
         \warp_checker_fence_regs_rd_cta_id[25><2] ,
         \warp_checker_fence_regs_rd_cta_id[25><1] ,
         \warp_checker_fence_regs_rd_cta_id[25><0] ,
         \warp_checker_fence_regs_rd_cta_id[24><3] ,
         \warp_checker_fence_regs_rd_cta_id[24><2] ,
         \warp_checker_fence_regs_rd_cta_id[24><1] ,
         \warp_checker_fence_regs_rd_cta_id[24><0] ,
         \warp_checker_fence_regs_rd_cta_id[23><3] ,
         \warp_checker_fence_regs_rd_cta_id[23><2] ,
         \warp_checker_fence_regs_rd_cta_id[23><1] ,
         \warp_checker_fence_regs_rd_cta_id[23><0] ,
         \warp_checker_fence_regs_rd_cta_id[22><3] ,
         \warp_checker_fence_regs_rd_cta_id[22><2] ,
         \warp_checker_fence_regs_rd_cta_id[22><1] ,
         \warp_checker_fence_regs_rd_cta_id[22><0] ,
         \warp_checker_fence_regs_rd_cta_id[21><3] ,
         \warp_checker_fence_regs_rd_cta_id[21><2] ,
         \warp_checker_fence_regs_rd_cta_id[21><1] ,
         \warp_checker_fence_regs_rd_cta_id[21><0] ,
         \warp_checker_fence_regs_rd_cta_id[20><3] ,
         \warp_checker_fence_regs_rd_cta_id[20><2] ,
         \warp_checker_fence_regs_rd_cta_id[20><1] ,
         \warp_checker_fence_regs_rd_cta_id[20><0] ,
         \warp_checker_fence_regs_rd_cta_id[19><3] ,
         \warp_checker_fence_regs_rd_cta_id[19><2] ,
         \warp_checker_fence_regs_rd_cta_id[19><1] ,
         \warp_checker_fence_regs_rd_cta_id[19><0] ,
         \warp_checker_fence_regs_rd_cta_id[18><3] ,
         \warp_checker_fence_regs_rd_cta_id[18><2] ,
         \warp_checker_fence_regs_rd_cta_id[18><1] ,
         \warp_checker_fence_regs_rd_cta_id[18><0] ,
         \warp_checker_fence_regs_rd_cta_id[17><3] ,
         \warp_checker_fence_regs_rd_cta_id[17><2] ,
         \warp_checker_fence_regs_rd_cta_id[17><1] ,
         \warp_checker_fence_regs_rd_cta_id[17><0] ,
         \warp_checker_fence_regs_rd_cta_id[16><3] ,
         \warp_checker_fence_regs_rd_cta_id[16><2] ,
         \warp_checker_fence_regs_rd_cta_id[16><1] ,
         \warp_checker_fence_regs_rd_cta_id[16><0] ,
         \warp_checker_fence_regs_rd_cta_id[15><3] ,
         \warp_checker_fence_regs_rd_cta_id[15><2] ,
         \warp_checker_fence_regs_rd_cta_id[15><1] ,
         \warp_checker_fence_regs_rd_cta_id[15><0] ,
         \warp_checker_fence_regs_rd_cta_id[14><3] ,
         \warp_checker_fence_regs_rd_cta_id[14><2] ,
         \warp_checker_fence_regs_rd_cta_id[14><1] ,
         \warp_checker_fence_regs_rd_cta_id[14><0] ,
         \warp_checker_fence_regs_rd_cta_id[13><3] ,
         \warp_checker_fence_regs_rd_cta_id[13><2] ,
         \warp_checker_fence_regs_rd_cta_id[13><1] ,
         \warp_checker_fence_regs_rd_cta_id[13><0] ,
         \warp_checker_fence_regs_rd_cta_id[12><3] ,
         \warp_checker_fence_regs_rd_cta_id[12><2] ,
         \warp_checker_fence_regs_rd_cta_id[12><1] ,
         \warp_checker_fence_regs_rd_cta_id[12><0] ,
         \warp_checker_fence_regs_rd_cta_id[11><3] ,
         \warp_checker_fence_regs_rd_cta_id[11><2] ,
         \warp_checker_fence_regs_rd_cta_id[11><1] ,
         \warp_checker_fence_regs_rd_cta_id[11><0] ,
         \warp_checker_fence_regs_rd_cta_id[10><3] ,
         \warp_checker_fence_regs_rd_cta_id[10><2] ,
         \warp_checker_fence_regs_rd_cta_id[10><1] ,
         \warp_checker_fence_regs_rd_cta_id[10><0] ,
         \warp_checker_fence_regs_rd_cta_id[9><3] ,
         \warp_checker_fence_regs_rd_cta_id[9><2] ,
         \warp_checker_fence_regs_rd_cta_id[9><1] ,
         \warp_checker_fence_regs_rd_cta_id[9><0] ,
         \warp_checker_fence_regs_rd_cta_id[8><3] ,
         \warp_checker_fence_regs_rd_cta_id[8><2] ,
         \warp_checker_fence_regs_rd_cta_id[8><1] ,
         \warp_checker_fence_regs_rd_cta_id[8><0] ,
         \warp_checker_fence_regs_rd_cta_id[7><3] ,
         \warp_checker_fence_regs_rd_cta_id[7><2] ,
         \warp_checker_fence_regs_rd_cta_id[7><1] ,
         \warp_checker_fence_regs_rd_cta_id[7><0] ,
         \warp_checker_fence_regs_rd_cta_id[6><3] ,
         \warp_checker_fence_regs_rd_cta_id[6><2] ,
         \warp_checker_fence_regs_rd_cta_id[6><1] ,
         \warp_checker_fence_regs_rd_cta_id[6><0] ,
         \warp_checker_fence_regs_rd_cta_id[5><3] ,
         \warp_checker_fence_regs_rd_cta_id[5><2] ,
         \warp_checker_fence_regs_rd_cta_id[5><1] ,
         \warp_checker_fence_regs_rd_cta_id[5><0] ,
         \warp_checker_fence_regs_rd_cta_id[4><3] ,
         \warp_checker_fence_regs_rd_cta_id[4><2] ,
         \warp_checker_fence_regs_rd_cta_id[4><1] ,
         \warp_checker_fence_regs_rd_cta_id[4><0] ,
         \warp_checker_fence_regs_rd_cta_id[3><3] ,
         \warp_checker_fence_regs_rd_cta_id[3><2] ,
         \warp_checker_fence_regs_rd_cta_id[3><1] ,
         \warp_checker_fence_regs_rd_cta_id[3><0] ,
         \warp_checker_fence_regs_rd_cta_id[2><3] ,
         \warp_checker_fence_regs_rd_cta_id[2><2] ,
         \warp_checker_fence_regs_rd_cta_id[2><1] ,
         \warp_checker_fence_regs_rd_cta_id[2><0] ,
         \warp_checker_fence_regs_rd_cta_id[1><3] ,
         \warp_checker_fence_regs_rd_cta_id[1><2] ,
         \warp_checker_fence_regs_rd_cta_id[1><1] ,
         \warp_checker_fence_regs_rd_cta_id[1><0] ,
         \warp_checker_fence_regs_rd_cta_id[0><3] ,
         \warp_checker_fence_regs_rd_cta_id[0><2] ,
         \warp_checker_fence_regs_rd_cta_id[0><1] ,
         \warp_checker_fence_regs_rd_cta_id[0><0] ,
         \fence_regs_rd_cta_id[31><3] , \fence_regs_rd_cta_id[31><2] ,
         \fence_regs_rd_cta_id[31><1] , \fence_regs_rd_cta_id[31><0] ,
         \fence_regs_rd_cta_id[30><3] , \fence_regs_rd_cta_id[30><2] ,
         \fence_regs_rd_cta_id[30><1] , \fence_regs_rd_cta_id[30><0] ,
         \fence_regs_rd_cta_id[29><3] , \fence_regs_rd_cta_id[29><2] ,
         \fence_regs_rd_cta_id[29><1] , \fence_regs_rd_cta_id[29><0] ,
         \fence_regs_rd_cta_id[28><3] , \fence_regs_rd_cta_id[28><2] ,
         \fence_regs_rd_cta_id[28><1] , \fence_regs_rd_cta_id[28><0] ,
         \fence_regs_rd_cta_id[27><3] , \fence_regs_rd_cta_id[27><2] ,
         \fence_regs_rd_cta_id[27><1] , \fence_regs_rd_cta_id[27><0] ,
         \fence_regs_rd_cta_id[26><3] , \fence_regs_rd_cta_id[26><2] ,
         \fence_regs_rd_cta_id[26><1] , \fence_regs_rd_cta_id[26><0] ,
         \fence_regs_rd_cta_id[25><3] , \fence_regs_rd_cta_id[25><2] ,
         \fence_regs_rd_cta_id[25><1] , \fence_regs_rd_cta_id[25><0] ,
         \fence_regs_rd_cta_id[24><3] , \fence_regs_rd_cta_id[24><2] ,
         \fence_regs_rd_cta_id[24><1] , \fence_regs_rd_cta_id[24><0] ,
         \fence_regs_rd_cta_id[23><3] , \fence_regs_rd_cta_id[23><2] ,
         \fence_regs_rd_cta_id[23><1] , \fence_regs_rd_cta_id[23><0] ,
         \fence_regs_rd_cta_id[22><3] , \fence_regs_rd_cta_id[22><2] ,
         \fence_regs_rd_cta_id[22><1] , \fence_regs_rd_cta_id[22><0] ,
         \fence_regs_rd_cta_id[21><3] , \fence_regs_rd_cta_id[21><2] ,
         \fence_regs_rd_cta_id[21><1] , \fence_regs_rd_cta_id[21><0] ,
         \fence_regs_rd_cta_id[20><3] , \fence_regs_rd_cta_id[20><2] ,
         \fence_regs_rd_cta_id[20><1] , \fence_regs_rd_cta_id[20><0] ,
         \fence_regs_rd_cta_id[19><3] , \fence_regs_rd_cta_id[19><2] ,
         \fence_regs_rd_cta_id[19><1] , \fence_regs_rd_cta_id[19><0] ,
         \fence_regs_rd_cta_id[18><3] , \fence_regs_rd_cta_id[18><2] ,
         \fence_regs_rd_cta_id[18><1] , \fence_regs_rd_cta_id[18><0] ,
         \fence_regs_rd_cta_id[17><3] , \fence_regs_rd_cta_id[17><2] ,
         \fence_regs_rd_cta_id[17><1] , \fence_regs_rd_cta_id[17><0] ,
         \fence_regs_rd_cta_id[16><3] , \fence_regs_rd_cta_id[16><2] ,
         \fence_regs_rd_cta_id[16><1] , \fence_regs_rd_cta_id[16><0] ,
         \fence_regs_rd_cta_id[15><3] , \fence_regs_rd_cta_id[15><2] ,
         \fence_regs_rd_cta_id[15><1] , \fence_regs_rd_cta_id[15><0] ,
         \fence_regs_rd_cta_id[14><3] , \fence_regs_rd_cta_id[14><2] ,
         \fence_regs_rd_cta_id[14><1] , \fence_regs_rd_cta_id[14><0] ,
         \fence_regs_rd_cta_id[13><3] , \fence_regs_rd_cta_id[13><2] ,
         \fence_regs_rd_cta_id[13><1] , \fence_regs_rd_cta_id[13><0] ,
         \fence_regs_rd_cta_id[12><3] , \fence_regs_rd_cta_id[12><2] ,
         \fence_regs_rd_cta_id[12><1] , \fence_regs_rd_cta_id[12><0] ,
         \fence_regs_rd_cta_id[11><3] , \fence_regs_rd_cta_id[11><2] ,
         \fence_regs_rd_cta_id[11><1] , \fence_regs_rd_cta_id[11><0] ,
         \fence_regs_rd_cta_id[10><3] , \fence_regs_rd_cta_id[10><2] ,
         \fence_regs_rd_cta_id[10><1] , \fence_regs_rd_cta_id[10><0] ,
         \fence_regs_rd_cta_id[9><3] , \fence_regs_rd_cta_id[9><2] ,
         \fence_regs_rd_cta_id[9><1] , \fence_regs_rd_cta_id[9><0] ,
         \fence_regs_rd_cta_id[8><3] , \fence_regs_rd_cta_id[8><2] ,
         \fence_regs_rd_cta_id[8><1] , \fence_regs_rd_cta_id[8><0] ,
         \fence_regs_rd_cta_id[7><3] , \fence_regs_rd_cta_id[7><2] ,
         \fence_regs_rd_cta_id[7><1] , \fence_regs_rd_cta_id[7><0] ,
         \fence_regs_rd_cta_id[6><3] , \fence_regs_rd_cta_id[6><2] ,
         \fence_regs_rd_cta_id[6><1] , \fence_regs_rd_cta_id[6><0] ,
         \fence_regs_rd_cta_id[5><3] , \fence_regs_rd_cta_id[5><2] ,
         \fence_regs_rd_cta_id[5><1] , \fence_regs_rd_cta_id[5><0] ,
         \fence_regs_rd_cta_id[4><3] , \fence_regs_rd_cta_id[4><2] ,
         \fence_regs_rd_cta_id[4><1] , \fence_regs_rd_cta_id[4><0] ,
         \fence_regs_rd_cta_id[3><3] , \fence_regs_rd_cta_id[3><2] ,
         \fence_regs_rd_cta_id[3><1] , \fence_regs_rd_cta_id[3><0] ,
         \fence_regs_rd_cta_id[2><3] , \fence_regs_rd_cta_id[2><2] ,
         \fence_regs_rd_cta_id[2><1] , \fence_regs_rd_cta_id[2><0] ,
         \fence_regs_rd_cta_id[1><3] , \fence_regs_rd_cta_id[1><2] ,
         \fence_regs_rd_cta_id[1><1] , \fence_regs_rd_cta_id[1><0] ,
         \fence_regs_rd_cta_id[0><3] , \fence_regs_rd_cta_id[0><2] ,
         \fence_regs_rd_cta_id[0><1] , \fence_regs_rd_cta_id[0><0] ,
         \fence_regs_wr_cta_id[31><3] , \fence_regs_wr_cta_id[31><2] ,
         \fence_regs_wr_cta_id[31><1] , \fence_regs_wr_cta_id[31><0] ,
         \fence_regs_wr_cta_id[30><3] , \fence_regs_wr_cta_id[30><2] ,
         \fence_regs_wr_cta_id[30><1] , \fence_regs_wr_cta_id[30><0] ,
         \fence_regs_wr_cta_id[29><3] , \fence_regs_wr_cta_id[29><2] ,
         \fence_regs_wr_cta_id[29><1] , \fence_regs_wr_cta_id[29><0] ,
         \fence_regs_wr_cta_id[28><3] , \fence_regs_wr_cta_id[28><2] ,
         \fence_regs_wr_cta_id[28><1] , \fence_regs_wr_cta_id[28><0] ,
         \fence_regs_wr_cta_id[27><3] , \fence_regs_wr_cta_id[27><2] ,
         \fence_regs_wr_cta_id[27><1] , \fence_regs_wr_cta_id[27><0] ,
         \fence_regs_wr_cta_id[26><3] , \fence_regs_wr_cta_id[26><2] ,
         \fence_regs_wr_cta_id[26><1] , \fence_regs_wr_cta_id[26><0] ,
         \fence_regs_wr_cta_id[25><3] , \fence_regs_wr_cta_id[25><2] ,
         \fence_regs_wr_cta_id[25><1] , \fence_regs_wr_cta_id[25><0] ,
         \fence_regs_wr_cta_id[24><3] , \fence_regs_wr_cta_id[24><2] ,
         \fence_regs_wr_cta_id[24><1] , \fence_regs_wr_cta_id[24><0] ,
         \fence_regs_wr_cta_id[23><3] , \fence_regs_wr_cta_id[23><2] ,
         \fence_regs_wr_cta_id[23><1] , \fence_regs_wr_cta_id[23><0] ,
         \fence_regs_wr_cta_id[22><3] , \fence_regs_wr_cta_id[22><2] ,
         \fence_regs_wr_cta_id[22><1] , \fence_regs_wr_cta_id[22><0] ,
         \fence_regs_wr_cta_id[21><3] , \fence_regs_wr_cta_id[21><2] ,
         \fence_regs_wr_cta_id[21><1] , \fence_regs_wr_cta_id[21><0] ,
         \fence_regs_wr_cta_id[20><3] , \fence_regs_wr_cta_id[20><2] ,
         \fence_regs_wr_cta_id[20><1] , \fence_regs_wr_cta_id[20><0] ,
         \fence_regs_wr_cta_id[19><3] , \fence_regs_wr_cta_id[19><2] ,
         \fence_regs_wr_cta_id[19><1] , \fence_regs_wr_cta_id[19><0] ,
         \fence_regs_wr_cta_id[18><3] , \fence_regs_wr_cta_id[18><2] ,
         \fence_regs_wr_cta_id[18><1] , \fence_regs_wr_cta_id[18><0] ,
         \fence_regs_wr_cta_id[17><3] , \fence_regs_wr_cta_id[17><2] ,
         \fence_regs_wr_cta_id[17><1] , \fence_regs_wr_cta_id[17><0] ,
         \fence_regs_wr_cta_id[16><3] , \fence_regs_wr_cta_id[16><2] ,
         \fence_regs_wr_cta_id[16><1] , \fence_regs_wr_cta_id[16><0] ,
         \fence_regs_wr_cta_id[15><3] , \fence_regs_wr_cta_id[15><2] ,
         \fence_regs_wr_cta_id[15><1] , \fence_regs_wr_cta_id[15><0] ,
         \fence_regs_wr_cta_id[14><3] , \fence_regs_wr_cta_id[14><2] ,
         \fence_regs_wr_cta_id[14><1] , \fence_regs_wr_cta_id[14><0] ,
         \fence_regs_wr_cta_id[13><3] , \fence_regs_wr_cta_id[13><2] ,
         \fence_regs_wr_cta_id[13><1] , \fence_regs_wr_cta_id[13><0] ,
         \fence_regs_wr_cta_id[12><3] , \fence_regs_wr_cta_id[12><2] ,
         \fence_regs_wr_cta_id[12><1] , \fence_regs_wr_cta_id[12><0] ,
         \fence_regs_wr_cta_id[11><3] , \fence_regs_wr_cta_id[11><2] ,
         \fence_regs_wr_cta_id[11><1] , \fence_regs_wr_cta_id[11><0] ,
         \fence_regs_wr_cta_id[10><3] , \fence_regs_wr_cta_id[10><2] ,
         \fence_regs_wr_cta_id[10><1] , \fence_regs_wr_cta_id[10><0] ,
         \fence_regs_wr_cta_id[9><3] , \fence_regs_wr_cta_id[9><2] ,
         \fence_regs_wr_cta_id[9><1] , \fence_regs_wr_cta_id[9><0] ,
         \fence_regs_wr_cta_id[8><3] , \fence_regs_wr_cta_id[8><2] ,
         \fence_regs_wr_cta_id[8><1] , \fence_regs_wr_cta_id[8><0] ,
         \fence_regs_wr_cta_id[7><3] , \fence_regs_wr_cta_id[7><2] ,
         \fence_regs_wr_cta_id[7><1] , \fence_regs_wr_cta_id[7><0] ,
         \fence_regs_wr_cta_id[6><3] , \fence_regs_wr_cta_id[6><2] ,
         \fence_regs_wr_cta_id[6><1] , \fence_regs_wr_cta_id[6><0] ,
         \fence_regs_wr_cta_id[5><3] , \fence_regs_wr_cta_id[5><2] ,
         \fence_regs_wr_cta_id[5><1] , \fence_regs_wr_cta_id[5><0] ,
         \fence_regs_wr_cta_id[4><3] , \fence_regs_wr_cta_id[4><2] ,
         \fence_regs_wr_cta_id[4><1] , \fence_regs_wr_cta_id[4><0] ,
         \fence_regs_wr_cta_id[3><3] , \fence_regs_wr_cta_id[3><2] ,
         \fence_regs_wr_cta_id[3><1] , \fence_regs_wr_cta_id[3><0] ,
         \fence_regs_wr_cta_id[2><3] , \fence_regs_wr_cta_id[2><2] ,
         \fence_regs_wr_cta_id[2><1] , \fence_regs_wr_cta_id[2><0] ,
         \fence_regs_wr_cta_id[1><3] , \fence_regs_wr_cta_id[1><2] ,
         \fence_regs_wr_cta_id[1><1] , \fence_regs_wr_cta_id[1><0] ,
         \fence_regs_wr_cta_id[0><3] , \fence_regs_wr_cta_id[0><2] ,
         \fence_regs_wr_cta_id[0><1] , \fence_regs_wr_cta_id[0><0] , n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n208, n211, n212, n213, n214, n215, n345, n346, n347, n348, n349,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n209, n210, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261;
  wire   [4:0] warp_gen_pool_addr;
  wire   [127:0] warp_gen_pool_wr_data;
  wire   [4:0] warp_gen_state_addr;
  wire   [31:0] warp_gen_fence_regs_cta_id_ld;
  wire   [31:0] warp_gen_fence_regs_fence_en_ld;
  wire   [31:0] warps_done_mask_int;
  wire   [4:0] warp_sched_pool_addr;
  wire   [4:0] warp_sched_state_addr;
  wire   [4:0] warp_pool_addr_b;
  wire   [127:0] warp_pool_wr_data_b;
  wire   [4:0] warp_state_addr_b;
  wire   [1:0] warp_state_wr_data_b;
  wire   [31:0] warp_checker_fence_regs_wr_fence_en;
  wire   [31:0] warp_checker_fence_regs_fence_en_ld;
  wire   [31:0] warp_checker_fence_regs_rd_fence_en;
  wire   [127:0] warp_pool_rd_data_a;
  wire   [1:0] warp_state_rd_data_a;
  wire   [31:0] fence_regs_rd_fence_en;
  wire   [31:0] fence_regs_cta_id_ld;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42;

  warp_generator uWarpGenerator ( .clk_in(clk_in), 
        .host_reset(n248), .en(warp_generator_en), .num_blocks_in(
        num_blocks_in), .warps_per_block_in(warps_per_block_in), 
        .shmem_base_addr_in(shared_mem_base_addr_in), .shmem_size_in(
        shared_mem_size_in), .gprs_size_in(gprs_size_in), .warp_pool_addr_out(
        warp_gen_pool_addr), .warp_pool_wr_en_out(warp_gen_pool_wr_en), 
        .warp_pool_wr_data_out({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, warp_gen_pool_wr_data[123:97], 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, warp_gen_pool_wr_data[63:0]}), 
        .warp_state_addr_out(warp_gen_state_addr), .warp_state_wr_en_out(
        warp_gen_state_wr_en), .fence_regs_cta_id_out({
        \warp_gen_fence_regs_wr_cta_id[31><3] , 
        \warp_gen_fence_regs_wr_cta_id[31><2] , 
        \warp_gen_fence_regs_wr_cta_id[31><1] , 
        \warp_gen_fence_regs_wr_cta_id[31><0] , 
        \warp_gen_fence_regs_wr_cta_id[30><3] , 
        \warp_gen_fence_regs_wr_cta_id[30><2] , 
        \warp_gen_fence_regs_wr_cta_id[30><1] , 
        \warp_gen_fence_regs_wr_cta_id[30><0] , 
        \warp_gen_fence_regs_wr_cta_id[29><3] , 
        \warp_gen_fence_regs_wr_cta_id[29><2] , 
        \warp_gen_fence_regs_wr_cta_id[29><1] , 
        \warp_gen_fence_regs_wr_cta_id[29><0] , 
        \warp_gen_fence_regs_wr_cta_id[28><3] , 
        \warp_gen_fence_regs_wr_cta_id[28><2] , 
        \warp_gen_fence_regs_wr_cta_id[28><1] , 
        \warp_gen_fence_regs_wr_cta_id[28><0] , 
        \warp_gen_fence_regs_wr_cta_id[27><3] , 
        \warp_gen_fence_regs_wr_cta_id[27><2] , 
        \warp_gen_fence_regs_wr_cta_id[27><1] , 
        \warp_gen_fence_regs_wr_cta_id[27><0] , 
        \warp_gen_fence_regs_wr_cta_id[26><3] , 
        \warp_gen_fence_regs_wr_cta_id[26><2] , 
        \warp_gen_fence_regs_wr_cta_id[26><1] , 
        \warp_gen_fence_regs_wr_cta_id[26><0] , 
        \warp_gen_fence_regs_wr_cta_id[25><3] , 
        \warp_gen_fence_regs_wr_cta_id[25><2] , 
        \warp_gen_fence_regs_wr_cta_id[25><1] , 
        \warp_gen_fence_regs_wr_cta_id[25><0] , 
        \warp_gen_fence_regs_wr_cta_id[24><3] , 
        \warp_gen_fence_regs_wr_cta_id[24><2] , 
        \warp_gen_fence_regs_wr_cta_id[24><1] , 
        \warp_gen_fence_regs_wr_cta_id[24><0] , 
        \warp_gen_fence_regs_wr_cta_id[23><3] , 
        \warp_gen_fence_regs_wr_cta_id[23><2] , 
        \warp_gen_fence_regs_wr_cta_id[23><1] , 
        \warp_gen_fence_regs_wr_cta_id[23><0] , 
        \warp_gen_fence_regs_wr_cta_id[22><3] , 
        \warp_gen_fence_regs_wr_cta_id[22><2] , 
        \warp_gen_fence_regs_wr_cta_id[22><1] , 
        \warp_gen_fence_regs_wr_cta_id[22><0] , 
        \warp_gen_fence_regs_wr_cta_id[21><3] , 
        \warp_gen_fence_regs_wr_cta_id[21><2] , 
        \warp_gen_fence_regs_wr_cta_id[21><1] , 
        \warp_gen_fence_regs_wr_cta_id[21><0] , 
        \warp_gen_fence_regs_wr_cta_id[20><3] , 
        \warp_gen_fence_regs_wr_cta_id[20><2] , 
        \warp_gen_fence_regs_wr_cta_id[20><1] , 
        \warp_gen_fence_regs_wr_cta_id[20><0] , 
        \warp_gen_fence_regs_wr_cta_id[19><3] , 
        \warp_gen_fence_regs_wr_cta_id[19><2] , 
        \warp_gen_fence_regs_wr_cta_id[19><1] , 
        \warp_gen_fence_regs_wr_cta_id[19><0] , 
        \warp_gen_fence_regs_wr_cta_id[18><3] , 
        \warp_gen_fence_regs_wr_cta_id[18><2] , 
        \warp_gen_fence_regs_wr_cta_id[18><1] , 
        \warp_gen_fence_regs_wr_cta_id[18><0] , 
        \warp_gen_fence_regs_wr_cta_id[17><3] , 
        \warp_gen_fence_regs_wr_cta_id[17><2] , 
        \warp_gen_fence_regs_wr_cta_id[17><1] , 
        \warp_gen_fence_regs_wr_cta_id[17><0] , 
        \warp_gen_fence_regs_wr_cta_id[16><3] , 
        \warp_gen_fence_regs_wr_cta_id[16><2] , 
        \warp_gen_fence_regs_wr_cta_id[16><1] , 
        \warp_gen_fence_regs_wr_cta_id[16><0] , 
        \warp_gen_fence_regs_wr_cta_id[15><3] , 
        \warp_gen_fence_regs_wr_cta_id[15><2] , 
        \warp_gen_fence_regs_wr_cta_id[15><1] , 
        \warp_gen_fence_regs_wr_cta_id[15><0] , 
        \warp_gen_fence_regs_wr_cta_id[14><3] , 
        \warp_gen_fence_regs_wr_cta_id[14><2] , 
        \warp_gen_fence_regs_wr_cta_id[14><1] , 
        \warp_gen_fence_regs_wr_cta_id[14><0] , 
        \warp_gen_fence_regs_wr_cta_id[13><3] , 
        \warp_gen_fence_regs_wr_cta_id[13><2] , 
        \warp_gen_fence_regs_wr_cta_id[13><1] , 
        \warp_gen_fence_regs_wr_cta_id[13><0] , 
        \warp_gen_fence_regs_wr_cta_id[12><3] , 
        \warp_gen_fence_regs_wr_cta_id[12><2] , 
        \warp_gen_fence_regs_wr_cta_id[12><1] , 
        \warp_gen_fence_regs_wr_cta_id[12><0] , 
        \warp_gen_fence_regs_wr_cta_id[11><3] , 
        \warp_gen_fence_regs_wr_cta_id[11><2] , 
        \warp_gen_fence_regs_wr_cta_id[11><1] , 
        \warp_gen_fence_regs_wr_cta_id[11><0] , 
        \warp_gen_fence_regs_wr_cta_id[10><3] , 
        \warp_gen_fence_regs_wr_cta_id[10><2] , 
        \warp_gen_fence_regs_wr_cta_id[10><1] , 
        \warp_gen_fence_regs_wr_cta_id[10><0] , 
        \warp_gen_fence_regs_wr_cta_id[9><3] , 
        \warp_gen_fence_regs_wr_cta_id[9><2] , 
        \warp_gen_fence_regs_wr_cta_id[9><1] , 
        \warp_gen_fence_regs_wr_cta_id[9><0] , 
        \warp_gen_fence_regs_wr_cta_id[8><3] , 
        \warp_gen_fence_regs_wr_cta_id[8><2] , 
        \warp_gen_fence_regs_wr_cta_id[8><1] , 
        \warp_gen_fence_regs_wr_cta_id[8><0] , 
        \warp_gen_fence_regs_wr_cta_id[7><3] , 
        \warp_gen_fence_regs_wr_cta_id[7><2] , 
        \warp_gen_fence_regs_wr_cta_id[7><1] , 
        \warp_gen_fence_regs_wr_cta_id[7><0] , 
        \warp_gen_fence_regs_wr_cta_id[6><3] , 
        \warp_gen_fence_regs_wr_cta_id[6><2] , 
        \warp_gen_fence_regs_wr_cta_id[6><1] , 
        \warp_gen_fence_regs_wr_cta_id[6><0] , 
        \warp_gen_fence_regs_wr_cta_id[5><3] , 
        \warp_gen_fence_regs_wr_cta_id[5><2] , 
        \warp_gen_fence_regs_wr_cta_id[5><1] , 
        \warp_gen_fence_regs_wr_cta_id[5><0] , 
        \warp_gen_fence_regs_wr_cta_id[4><3] , 
        \warp_gen_fence_regs_wr_cta_id[4><2] , 
        \warp_gen_fence_regs_wr_cta_id[4><1] , 
        \warp_gen_fence_regs_wr_cta_id[4><0] , 
        \warp_gen_fence_regs_wr_cta_id[3><3] , 
        \warp_gen_fence_regs_wr_cta_id[3><2] , 
        \warp_gen_fence_regs_wr_cta_id[3><1] , 
        \warp_gen_fence_regs_wr_cta_id[3><0] , 
        \warp_gen_fence_regs_wr_cta_id[2><3] , 
        \warp_gen_fence_regs_wr_cta_id[2><2] , 
        \warp_gen_fence_regs_wr_cta_id[2><1] , 
        \warp_gen_fence_regs_wr_cta_id[2><0] , 
        \warp_gen_fence_regs_wr_cta_id[1><3] , 
        \warp_gen_fence_regs_wr_cta_id[1><2] , 
        \warp_gen_fence_regs_wr_cta_id[1><1] , 
        \warp_gen_fence_regs_wr_cta_id[1><0] , 
        \warp_gen_fence_regs_wr_cta_id[0><3] , 
        \warp_gen_fence_regs_wr_cta_id[0><2] , 
        \warp_gen_fence_regs_wr_cta_id[0><1] , 
        \warp_gen_fence_regs_wr_cta_id[0><0] }), .fence_regs_cta_id_ld(
        warp_gen_fence_regs_cta_id_ld), .fence_regs_fence_en_ld(
        warp_gen_fence_regs_fence_en_ld), .num_warps_out(num_warps_out), 
        .warp_gen_done(warp_generator_done) );
		
  warp_scheduler uWarpScheduler ( .clk_in(clk_in), 
        .host_reset(n248), .reset(n164), .pipeline_stall_in(pipeline_stall_in), 
        .num_blocks_in(num_blocks_in), .num_warps_in(num_warps_out), 
        .gprs_size_in(gprs_size_in), .warps_done_mask_in(warps_done_mask_int), 
        .warp_pool_addr_out(warp_sched_pool_addr), .warp_pool_rd_data_in(
        warp_pool_rd_data_a), .warp_state_addr_out(warp_sched_state_addr), 
        .warp_state_wr_en_out(warp_sched_state_wr_en), 
        .warp_state_wr_data_out({SYNOPSYS_UNCONNECTED__37, 
        \warp_sched_state_wr_data[0] }), .warp_state_rd_data_in(
        warp_state_rd_data_a), .program_cntr_out(program_cntr_out), 
        .warp_id_out(warp_id_out), .warp_lane_id_out(warp_lane_id_out), 
        .cta_id_out(cta_id_out), .initial_mask_out(initial_mask_out), 
        .current_mask_out(current_mask_out), .shmem_base_addr_out(
        shmem_base_addr_out), .gprs_size_out(gprs_size_out), 
        .gprs_base_addr_out(gprs_base_addr_out), .done(warp_scheduler_done), 
        .pipeline_warpunit_done(pipeline_warpunit_done), .fetch_en(fetch_en)
         );
  warp_checker uWarpChecker ( .clk_in(clk_in), .host_reset(
        n249), .reset(n164), .en(pipeline_write_done), .warp_id_in(warp_id_in), 
        .warp_lane_id_in(warp_lane_id_in), .cta_id_in(cta_id_in), 
        .initial_mask_in(initial_mask_in), .current_mask_in(current_mask_in), 
        .shmem_base_addr_in(shmem_base_addr_in), .gprs_base_addr_in(
        gprs_base_addr_in), .next_pc_in(next_pc_in), .warp_state_in(
        warp_state_in), .warps_per_block_in(warps_per_block_in), 
        .warp_pool_addr_out(warp_pool_addr_b), .warp_pool_wr_en_out(
        warp_pool_wr_en_b), .warp_pool_wr_data_out({SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, warp_pool_wr_data_b[123:97], 
        SYNOPSYS_UNCONNECTED__42, warp_pool_wr_data_b[95:0]}), 
        .warp_state_addr_out(warp_state_addr_b), .warp_state_wr_en_out(
        warp_state_wr_en_b), .warp_state_wr_data_out(warp_state_wr_data_b), 
        .fence_regs_fence_en_out(warp_checker_fence_regs_wr_fence_en), 
        .fence_regs_fence_en_ld(warp_checker_fence_regs_fence_en_ld), 
        .fence_regs_cta_id_in({\warp_checker_fence_regs_rd_cta_id[31><3] , 
        \warp_checker_fence_regs_rd_cta_id[31><2] , 
        \warp_checker_fence_regs_rd_cta_id[31><1] , 
        \warp_checker_fence_regs_rd_cta_id[31><0] , 
        \warp_checker_fence_regs_rd_cta_id[30><3] , 
        \warp_checker_fence_regs_rd_cta_id[30><2] , 
        \warp_checker_fence_regs_rd_cta_id[30><1] , 
        \warp_checker_fence_regs_rd_cta_id[30><0] , 
        \warp_checker_fence_regs_rd_cta_id[29><3] , 
        \warp_checker_fence_regs_rd_cta_id[29><2] , 
        \warp_checker_fence_regs_rd_cta_id[29><1] , 
        \warp_checker_fence_regs_rd_cta_id[29><0] , 
        \warp_checker_fence_regs_rd_cta_id[28><3] , 
        \warp_checker_fence_regs_rd_cta_id[28><2] , 
        \warp_checker_fence_regs_rd_cta_id[28><1] , 
        \warp_checker_fence_regs_rd_cta_id[28><0] , 
        \warp_checker_fence_regs_rd_cta_id[27><3] , 
        \warp_checker_fence_regs_rd_cta_id[27><2] , 
        \warp_checker_fence_regs_rd_cta_id[27><1] , 
        \warp_checker_fence_regs_rd_cta_id[27><0] , 
        \warp_checker_fence_regs_rd_cta_id[26><3] , 
        \warp_checker_fence_regs_rd_cta_id[26><2] , 
        \warp_checker_fence_regs_rd_cta_id[26><1] , 
        \warp_checker_fence_regs_rd_cta_id[26><0] , 
        \warp_checker_fence_regs_rd_cta_id[25><3] , 
        \warp_checker_fence_regs_rd_cta_id[25><2] , 
        \warp_checker_fence_regs_rd_cta_id[25><1] , 
        \warp_checker_fence_regs_rd_cta_id[25><0] , 
        \warp_checker_fence_regs_rd_cta_id[24><3] , 
        \warp_checker_fence_regs_rd_cta_id[24><2] , 
        \warp_checker_fence_regs_rd_cta_id[24><1] , 
        \warp_checker_fence_regs_rd_cta_id[24><0] , 
        \warp_checker_fence_regs_rd_cta_id[23><3] , 
        \warp_checker_fence_regs_rd_cta_id[23><2] , 
        \warp_checker_fence_regs_rd_cta_id[23><1] , 
        \warp_checker_fence_regs_rd_cta_id[23><0] , 
        \warp_checker_fence_regs_rd_cta_id[22><3] , 
        \warp_checker_fence_regs_rd_cta_id[22><2] , 
        \warp_checker_fence_regs_rd_cta_id[22><1] , 
        \warp_checker_fence_regs_rd_cta_id[22><0] , 
        \warp_checker_fence_regs_rd_cta_id[21><3] , 
        \warp_checker_fence_regs_rd_cta_id[21><2] , 
        \warp_checker_fence_regs_rd_cta_id[21><1] , 
        \warp_checker_fence_regs_rd_cta_id[21><0] , 
        \warp_checker_fence_regs_rd_cta_id[20><3] , 
        \warp_checker_fence_regs_rd_cta_id[20><2] , 
        \warp_checker_fence_regs_rd_cta_id[20><1] , 
        \warp_checker_fence_regs_rd_cta_id[20><0] , 
        \warp_checker_fence_regs_rd_cta_id[19><3] , 
        \warp_checker_fence_regs_rd_cta_id[19><2] , 
        \warp_checker_fence_regs_rd_cta_id[19><1] , 
        \warp_checker_fence_regs_rd_cta_id[19><0] , 
        \warp_checker_fence_regs_rd_cta_id[18><3] , 
        \warp_checker_fence_regs_rd_cta_id[18><2] , 
        \warp_checker_fence_regs_rd_cta_id[18><1] , 
        \warp_checker_fence_regs_rd_cta_id[18><0] , 
        \warp_checker_fence_regs_rd_cta_id[17><3] , 
        \warp_checker_fence_regs_rd_cta_id[17><2] , 
        \warp_checker_fence_regs_rd_cta_id[17><1] , 
        \warp_checker_fence_regs_rd_cta_id[17><0] , 
        \warp_checker_fence_regs_rd_cta_id[16><3] , 
        \warp_checker_fence_regs_rd_cta_id[16><2] , 
        \warp_checker_fence_regs_rd_cta_id[16><1] , 
        \warp_checker_fence_regs_rd_cta_id[16><0] , 
        \warp_checker_fence_regs_rd_cta_id[15><3] , 
        \warp_checker_fence_regs_rd_cta_id[15><2] , 
        \warp_checker_fence_regs_rd_cta_id[15><1] , 
        \warp_checker_fence_regs_rd_cta_id[15><0] , 
        \warp_checker_fence_regs_rd_cta_id[14><3] , 
        \warp_checker_fence_regs_rd_cta_id[14><2] , 
        \warp_checker_fence_regs_rd_cta_id[14><1] , 
        \warp_checker_fence_regs_rd_cta_id[14><0] , 
        \warp_checker_fence_regs_rd_cta_id[13><3] , 
        \warp_checker_fence_regs_rd_cta_id[13><2] , 
        \warp_checker_fence_regs_rd_cta_id[13><1] , 
        \warp_checker_fence_regs_rd_cta_id[13><0] , 
        \warp_checker_fence_regs_rd_cta_id[12><3] , 
        \warp_checker_fence_regs_rd_cta_id[12><2] , 
        \warp_checker_fence_regs_rd_cta_id[12><1] , 
        \warp_checker_fence_regs_rd_cta_id[12><0] , 
        \warp_checker_fence_regs_rd_cta_id[11><3] , 
        \warp_checker_fence_regs_rd_cta_id[11><2] , 
        \warp_checker_fence_regs_rd_cta_id[11><1] , 
        \warp_checker_fence_regs_rd_cta_id[11><0] , 
        \warp_checker_fence_regs_rd_cta_id[10><3] , 
        \warp_checker_fence_regs_rd_cta_id[10><2] , 
        \warp_checker_fence_regs_rd_cta_id[10><1] , 
        \warp_checker_fence_regs_rd_cta_id[10><0] , 
        \warp_checker_fence_regs_rd_cta_id[9><3] , 
        \warp_checker_fence_regs_rd_cta_id[9><2] , 
        \warp_checker_fence_regs_rd_cta_id[9><1] , 
        \warp_checker_fence_regs_rd_cta_id[9><0] , 
        \warp_checker_fence_regs_rd_cta_id[8><3] , 
        \warp_checker_fence_regs_rd_cta_id[8><2] , 
        \warp_checker_fence_regs_rd_cta_id[8><1] , 
        \warp_checker_fence_regs_rd_cta_id[8><0] , 
        \warp_checker_fence_regs_rd_cta_id[7><3] , 
        \warp_checker_fence_regs_rd_cta_id[7><2] , 
        \warp_checker_fence_regs_rd_cta_id[7><1] , 
        \warp_checker_fence_regs_rd_cta_id[7><0] , 
        \warp_checker_fence_regs_rd_cta_id[6><3] , 
        \warp_checker_fence_regs_rd_cta_id[6><2] , 
        \warp_checker_fence_regs_rd_cta_id[6><1] , 
        \warp_checker_fence_regs_rd_cta_id[6><0] , 
        \warp_checker_fence_regs_rd_cta_id[5><3] , 
        \warp_checker_fence_regs_rd_cta_id[5><2] , 
        \warp_checker_fence_regs_rd_cta_id[5><1] , 
        \warp_checker_fence_regs_rd_cta_id[5><0] , 
        \warp_checker_fence_regs_rd_cta_id[4><3] , 
        \warp_checker_fence_regs_rd_cta_id[4><2] , 
        \warp_checker_fence_regs_rd_cta_id[4><1] , 
        \warp_checker_fence_regs_rd_cta_id[4><0] , 
        \warp_checker_fence_regs_rd_cta_id[3><3] , 
        \warp_checker_fence_regs_rd_cta_id[3><2] , 
        \warp_checker_fence_regs_rd_cta_id[3><1] , 
        \warp_checker_fence_regs_rd_cta_id[3><0] , 
        \warp_checker_fence_regs_rd_cta_id[2><3] , 
        \warp_checker_fence_regs_rd_cta_id[2><2] , 
        \warp_checker_fence_regs_rd_cta_id[2><1] , 
        \warp_checker_fence_regs_rd_cta_id[2><0] , 
        \warp_checker_fence_regs_rd_cta_id[1><3] , 
        \warp_checker_fence_regs_rd_cta_id[1><2] , 
        \warp_checker_fence_regs_rd_cta_id[1><1] , 
        \warp_checker_fence_regs_rd_cta_id[1><0] , 
        \warp_checker_fence_regs_rd_cta_id[0><3] , 
        \warp_checker_fence_regs_rd_cta_id[0><2] , 
        \warp_checker_fence_regs_rd_cta_id[0><1] , 
        \warp_checker_fence_regs_rd_cta_id[0><0] }), .fence_regs_fence_en_in(
        warp_checker_fence_regs_rd_fence_en), .warps_done_mask_out(
        warps_done_mask_int), .pipeline_stall_out(pipeline_stall_out) );
  dp_regfile_RAM_SIZE32_RAM_A_WIDTH5_RAM_D_WIDTH128_1 uWarpPoolMemory ( .clk(
        clk_in), .rst(n249), .addr_a({n259, n253, n255, n261, n257}), .din_a({
        1'b0, 1'b0, 1'b0, 1'b0, n88, n87, n86, n85, n84, n83, n82, n80, n79, 
        n78, n77, n76, n75, n74, n73, n72, n71, n70, n69, n68, n67, n66, n65, 
        n152, n151, n150, n149, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, n148, n147, n146, n145, n144, n143, n142, n141, n140, n139, n138, 
        n137, n104, n103, n102, n101, n100, n99, n98, n97, n96, n95, n94, n93, 
        n92, n91, n90, n136, n135, n134, n133, n132, n131, n130, n129, n128, 
        n127, n126, n125, n124, n123, n122, n121, n120, n119, n118, n117, n116, 
        n115, n114, n113, n112, n111, n110, n109, n108, n107, n106, n105, n156, 
        n155, n154, n153, n81}), .we_a(n89), .addr_b(warp_pool_addr_b), 
        .din_b({1'b0, 1'b0, 1'b0, 1'b0, warp_pool_wr_data_b[123:97], 1'b0, 
        warp_pool_wr_data_b[95:0]}), .we_b(warp_pool_wr_en_b), .dout_a(
        warp_pool_rd_data_a) );
  dp_regfile_RAM_SIZE32_RAM_A_WIDTH5_RAM_D_WIDTH2_1 uWarpStateMemory ( .clk(
        clk_in), .rst(n249), .addr_a({n258, n252, n254, n260, n256}), .din_a({
        1'b0, n157}), .we_a(n251), .addr_b(warp_state_addr_b), .din_b(
        warp_state_wr_data_b), .we_b(warp_state_wr_en_b), .dout_a(
        warp_state_rd_data_a) );
  fence_registers_1_0 uFenceRegisters_0 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[0><3] , \fence_regs_wr_cta_id[0><2] , 
        \fence_regs_wr_cta_id[0><1] , \fence_regs_wr_cta_id[0><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[0]), .fence_en_in(n55), .fence_en_ld(
        n1), .cta_id_out({\fence_regs_rd_cta_id[0><3] , 
        \fence_regs_rd_cta_id[0><2] , \fence_regs_rd_cta_id[0><1] , 
        \fence_regs_rd_cta_id[0><0] }), .fence_en_out(
        fence_regs_rd_fence_en[0]) );
  fence_registers_1_31 uFenceRegisters_1 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[1><3] , \fence_regs_wr_cta_id[1><2] , 
        \fence_regs_wr_cta_id[1><1] , \fence_regs_wr_cta_id[1><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[1]), .fence_en_in(n33), .fence_en_ld(
        n2), .cta_id_out({\fence_regs_rd_cta_id[1><3] , 
        \fence_regs_rd_cta_id[1><2] , \fence_regs_rd_cta_id[1><1] , 
        \fence_regs_rd_cta_id[1><0] }), .fence_en_out(
        fence_regs_rd_fence_en[1]) );
  fence_registers_1_30 uFenceRegisters_2 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[2><3] , \fence_regs_wr_cta_id[2><2] , 
        \fence_regs_wr_cta_id[2><1] , \fence_regs_wr_cta_id[2><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[2]), .fence_en_in(n34), .fence_en_ld(
        n3), .cta_id_out({\fence_regs_rd_cta_id[2><3] , 
        \fence_regs_rd_cta_id[2><2] , \fence_regs_rd_cta_id[2><1] , 
        \fence_regs_rd_cta_id[2><0] }), .fence_en_out(
        fence_regs_rd_fence_en[2]) );
  fence_registers_1_29 uFenceRegisters_3 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[3><3] , \fence_regs_wr_cta_id[3><2] , 
        \fence_regs_wr_cta_id[3><1] , \fence_regs_wr_cta_id[3><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[3]), .fence_en_in(n56), .fence_en_ld(
        n4), .cta_id_out({\fence_regs_rd_cta_id[3><3] , 
        \fence_regs_rd_cta_id[3><2] , \fence_regs_rd_cta_id[3><1] , 
        \fence_regs_rd_cta_id[3><0] }), .fence_en_out(
        fence_regs_rd_fence_en[3]) );
  fence_registers_1_28 uFenceRegisters_4 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[4><3] , \fence_regs_wr_cta_id[4><2] , 
        \fence_regs_wr_cta_id[4><1] , \fence_regs_wr_cta_id[4><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[4]), .fence_en_in(n35), .fence_en_ld(
        n5), .cta_id_out({\fence_regs_rd_cta_id[4><3] , 
        \fence_regs_rd_cta_id[4><2] , \fence_regs_rd_cta_id[4><1] , 
        \fence_regs_rd_cta_id[4><0] }), .fence_en_out(
        fence_regs_rd_fence_en[4]) );
  fence_registers_1_27 uFenceRegisters_5 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[5><3] , \fence_regs_wr_cta_id[5><2] , 
        \fence_regs_wr_cta_id[5><1] , \fence_regs_wr_cta_id[5><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[5]), .fence_en_in(n36), .fence_en_ld(
        n6), .cta_id_out({\fence_regs_rd_cta_id[5><3] , 
        \fence_regs_rd_cta_id[5><2] , \fence_regs_rd_cta_id[5><1] , 
        \fence_regs_rd_cta_id[5><0] }), .fence_en_out(
        fence_regs_rd_fence_en[5]) );
  fence_registers_1_26 uFenceRegisters_6 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[6><3] , \fence_regs_wr_cta_id[6><2] , 
        \fence_regs_wr_cta_id[6><1] , \fence_regs_wr_cta_id[6><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[6]), .fence_en_in(n37), .fence_en_ld(
        n7), .cta_id_out({\fence_regs_rd_cta_id[6><3] , 
        \fence_regs_rd_cta_id[6><2] , \fence_regs_rd_cta_id[6><1] , 
        \fence_regs_rd_cta_id[6><0] }), .fence_en_out(
        fence_regs_rd_fence_en[6]) );
  fence_registers_1_25 uFenceRegisters_7 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[7><3] , \fence_regs_wr_cta_id[7><2] , 
        \fence_regs_wr_cta_id[7><1] , \fence_regs_wr_cta_id[7><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[7]), .fence_en_in(n38), .fence_en_ld(
        n8), .cta_id_out({\fence_regs_rd_cta_id[7><3] , 
        \fence_regs_rd_cta_id[7><2] , \fence_regs_rd_cta_id[7><1] , 
        \fence_regs_rd_cta_id[7><0] }), .fence_en_out(
        fence_regs_rd_fence_en[7]) );
  fence_registers_1_24 uFenceRegisters_8 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[8><3] , \fence_regs_wr_cta_id[8><2] , 
        \fence_regs_wr_cta_id[8><1] , \fence_regs_wr_cta_id[8><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[8]), .fence_en_in(n39), .fence_en_ld(
        n9), .cta_id_out({\fence_regs_rd_cta_id[8><3] , 
        \fence_regs_rd_cta_id[8><2] , \fence_regs_rd_cta_id[8><1] , 
        \fence_regs_rd_cta_id[8><0] }), .fence_en_out(
        fence_regs_rd_fence_en[8]) );
  fence_registers_1_23 uFenceRegisters_9 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[9><3] , \fence_regs_wr_cta_id[9><2] , 
        \fence_regs_wr_cta_id[9><1] , \fence_regs_wr_cta_id[9><0] }), 
        .cta_id_ld(fence_regs_cta_id_ld[9]), .fence_en_in(n57), .fence_en_ld(
        n10), .cta_id_out({\fence_regs_rd_cta_id[9><3] , 
        \fence_regs_rd_cta_id[9><2] , \fence_regs_rd_cta_id[9><1] , 
        \fence_regs_rd_cta_id[9><0] }), .fence_en_out(
        fence_regs_rd_fence_en[9]) );
  fence_registers_1_22 uFenceRegisters_10 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[10><3] , 
        \fence_regs_wr_cta_id[10><2] , \fence_regs_wr_cta_id[10><1] , 
        \fence_regs_wr_cta_id[10><0] }), .cta_id_ld(fence_regs_cta_id_ld[10]), 
        .fence_en_in(n40), .fence_en_ld(n11), .cta_id_out({
        \fence_regs_rd_cta_id[10><3] , \fence_regs_rd_cta_id[10><2] , 
        \fence_regs_rd_cta_id[10><1] , \fence_regs_rd_cta_id[10><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[10]) );
  fence_registers_1_21 uFenceRegisters_11 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[11><3] , 
        \fence_regs_wr_cta_id[11><2] , \fence_regs_wr_cta_id[11><1] , 
        \fence_regs_wr_cta_id[11><0] }), .cta_id_ld(fence_regs_cta_id_ld[11]), 
        .fence_en_in(n41), .fence_en_ld(n12), .cta_id_out({
        \fence_regs_rd_cta_id[11><3] , \fence_regs_rd_cta_id[11><2] , 
        \fence_regs_rd_cta_id[11><1] , \fence_regs_rd_cta_id[11><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[11]) );
  fence_registers_1_20 uFenceRegisters_12 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[12><3] , 
        \fence_regs_wr_cta_id[12><2] , \fence_regs_wr_cta_id[12><1] , 
        \fence_regs_wr_cta_id[12><0] }), .cta_id_ld(fence_regs_cta_id_ld[12]), 
        .fence_en_in(n62), .fence_en_ld(n13), .cta_id_out({
        \fence_regs_rd_cta_id[12><3] , \fence_regs_rd_cta_id[12><2] , 
        \fence_regs_rd_cta_id[12><1] , \fence_regs_rd_cta_id[12><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[12]) );
  fence_registers_1_19 uFenceRegisters_13 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[13><3] , 
        \fence_regs_wr_cta_id[13><2] , \fence_regs_wr_cta_id[13><1] , 
        \fence_regs_wr_cta_id[13><0] }), .cta_id_ld(fence_regs_cta_id_ld[13]), 
        .fence_en_in(n42), .fence_en_ld(n14), .cta_id_out({
        \fence_regs_rd_cta_id[13><3] , \fence_regs_rd_cta_id[13><2] , 
        \fence_regs_rd_cta_id[13><1] , \fence_regs_rd_cta_id[13><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[13]) );
  fence_registers_1_18 uFenceRegisters_14 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[14><3] , 
        \fence_regs_wr_cta_id[14><2] , \fence_regs_wr_cta_id[14><1] , 
        \fence_regs_wr_cta_id[14><0] }), .cta_id_ld(fence_regs_cta_id_ld[14]), 
        .fence_en_in(n43), .fence_en_ld(n15), .cta_id_out({
        \fence_regs_rd_cta_id[14><3] , \fence_regs_rd_cta_id[14><2] , 
        \fence_regs_rd_cta_id[14><1] , \fence_regs_rd_cta_id[14><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[14]) );
  fence_registers_1_17 uFenceRegisters_15 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[15><3] , 
        \fence_regs_wr_cta_id[15><2] , \fence_regs_wr_cta_id[15><1] , 
        \fence_regs_wr_cta_id[15><0] }), .cta_id_ld(fence_regs_cta_id_ld[15]), 
        .fence_en_in(n58), .fence_en_ld(n16), .cta_id_out({
        \fence_regs_rd_cta_id[15><3] , \fence_regs_rd_cta_id[15><2] , 
        \fence_regs_rd_cta_id[15><1] , \fence_regs_rd_cta_id[15><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[15]) );
  fence_registers_1_16 uFenceRegisters_16 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[16><3] , 
        \fence_regs_wr_cta_id[16><2] , \fence_regs_wr_cta_id[16><1] , 
        \fence_regs_wr_cta_id[16><0] }), .cta_id_ld(fence_regs_cta_id_ld[16]), 
        .fence_en_in(n44), .fence_en_ld(n17), .cta_id_out({
        \fence_regs_rd_cta_id[16><3] , \fence_regs_rd_cta_id[16><2] , 
        \fence_regs_rd_cta_id[16><1] , \fence_regs_rd_cta_id[16><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[16]) );
  fence_registers_1_15 uFenceRegisters_17 ( .clk_in(clk_in), .host_reset(n249), 
        .cta_id_in({\fence_regs_wr_cta_id[17><3] , 
        \fence_regs_wr_cta_id[17><2] , \fence_regs_wr_cta_id[17><1] , 
        \fence_regs_wr_cta_id[17><0] }), .cta_id_ld(fence_regs_cta_id_ld[17]), 
        .fence_en_in(n63), .fence_en_ld(n18), .cta_id_out({
        \fence_regs_rd_cta_id[17><3] , \fence_regs_rd_cta_id[17><2] , 
        \fence_regs_rd_cta_id[17><1] , \fence_regs_rd_cta_id[17><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[17]) );
  fence_registers_1_14 uFenceRegisters_18 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[18><3] , 
        \fence_regs_wr_cta_id[18><2] , \fence_regs_wr_cta_id[18><1] , 
        \fence_regs_wr_cta_id[18><0] }), .cta_id_ld(fence_regs_cta_id_ld[18]), 
        .fence_en_in(n45), .fence_en_ld(n19), .cta_id_out({
        \fence_regs_rd_cta_id[18><3] , \fence_regs_rd_cta_id[18><2] , 
        \fence_regs_rd_cta_id[18><1] , \fence_regs_rd_cta_id[18><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[18]) );
  fence_registers_1_13 uFenceRegisters_19 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[19><3] , 
        \fence_regs_wr_cta_id[19><2] , \fence_regs_wr_cta_id[19><1] , 
        \fence_regs_wr_cta_id[19><0] }), .cta_id_ld(fence_regs_cta_id_ld[19]), 
        .fence_en_in(n46), .fence_en_ld(n20), .cta_id_out({
        \fence_regs_rd_cta_id[19><3] , \fence_regs_rd_cta_id[19><2] , 
        \fence_regs_rd_cta_id[19><1] , \fence_regs_rd_cta_id[19><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[19]) );
  fence_registers_1_12 uFenceRegisters_20 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[20><3] , 
        \fence_regs_wr_cta_id[20><2] , \fence_regs_wr_cta_id[20><1] , 
        \fence_regs_wr_cta_id[20><0] }), .cta_id_ld(fence_regs_cta_id_ld[20]), 
        .fence_en_in(n47), .fence_en_ld(n21), .cta_id_out({
        \fence_regs_rd_cta_id[20><3] , \fence_regs_rd_cta_id[20><2] , 
        \fence_regs_rd_cta_id[20><1] , \fence_regs_rd_cta_id[20><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[20]) );
  fence_registers_1_11 uFenceRegisters_21 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[21><3] , 
        \fence_regs_wr_cta_id[21><2] , \fence_regs_wr_cta_id[21><1] , 
        \fence_regs_wr_cta_id[21><0] }), .cta_id_ld(fence_regs_cta_id_ld[21]), 
        .fence_en_in(n48), .fence_en_ld(n22), .cta_id_out({
        \fence_regs_rd_cta_id[21><3] , \fence_regs_rd_cta_id[21><2] , 
        \fence_regs_rd_cta_id[21><1] , \fence_regs_rd_cta_id[21><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[21]) );
  fence_registers_1_10 uFenceRegisters_22 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[22><3] , 
        \fence_regs_wr_cta_id[22><2] , \fence_regs_wr_cta_id[22><1] , 
        \fence_regs_wr_cta_id[22><0] }), .cta_id_ld(fence_regs_cta_id_ld[22]), 
        .fence_en_in(n49), .fence_en_ld(n23), .cta_id_out({
        \fence_regs_rd_cta_id[22><3] , \fence_regs_rd_cta_id[22><2] , 
        \fence_regs_rd_cta_id[22><1] , \fence_regs_rd_cta_id[22><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[22]) );
  fence_registers_1_9 uFenceRegisters_23 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[23><3] , 
        \fence_regs_wr_cta_id[23><2] , \fence_regs_wr_cta_id[23><1] , 
        \fence_regs_wr_cta_id[23><0] }), .cta_id_ld(fence_regs_cta_id_ld[23]), 
        .fence_en_in(n50), .fence_en_ld(n24), .cta_id_out({
        \fence_regs_rd_cta_id[23><3] , \fence_regs_rd_cta_id[23><2] , 
        \fence_regs_rd_cta_id[23><1] , \fence_regs_rd_cta_id[23><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[23]) );
  fence_registers_1_8 uFenceRegisters_24 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[24><3] , 
        \fence_regs_wr_cta_id[24><2] , \fence_regs_wr_cta_id[24><1] , 
        \fence_regs_wr_cta_id[24><0] }), .cta_id_ld(fence_regs_cta_id_ld[24]), 
        .fence_en_in(n51), .fence_en_ld(n25), .cta_id_out({
        \fence_regs_rd_cta_id[24><3] , \fence_regs_rd_cta_id[24><2] , 
        \fence_regs_rd_cta_id[24><1] , \fence_regs_rd_cta_id[24><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[24]) );
  fence_registers_1_7 uFenceRegisters_25 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[25><3] , 
        \fence_regs_wr_cta_id[25><2] , \fence_regs_wr_cta_id[25><1] , 
        \fence_regs_wr_cta_id[25><0] }), .cta_id_ld(fence_regs_cta_id_ld[25]), 
        .fence_en_in(n52), .fence_en_ld(n26), .cta_id_out({
        \fence_regs_rd_cta_id[25><3] , \fence_regs_rd_cta_id[25><2] , 
        \fence_regs_rd_cta_id[25><1] , \fence_regs_rd_cta_id[25><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[25]) );
  fence_registers_1_6 uFenceRegisters_26 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[26><3] , 
        \fence_regs_wr_cta_id[26><2] , \fence_regs_wr_cta_id[26><1] , 
        \fence_regs_wr_cta_id[26><0] }), .cta_id_ld(fence_regs_cta_id_ld[26]), 
        .fence_en_in(n53), .fence_en_ld(n27), .cta_id_out({
        \fence_regs_rd_cta_id[26><3] , \fence_regs_rd_cta_id[26><2] , 
        \fence_regs_rd_cta_id[26><1] , \fence_regs_rd_cta_id[26><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[26]) );
  fence_registers_1_5 uFenceRegisters_27 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[27><3] , 
        \fence_regs_wr_cta_id[27><2] , \fence_regs_wr_cta_id[27><1] , 
        \fence_regs_wr_cta_id[27><0] }), .cta_id_ld(fence_regs_cta_id_ld[27]), 
        .fence_en_in(n54), .fence_en_ld(n28), .cta_id_out({
        \fence_regs_rd_cta_id[27><3] , \fence_regs_rd_cta_id[27><2] , 
        \fence_regs_rd_cta_id[27><1] , \fence_regs_rd_cta_id[27><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[27]) );
  fence_registers_1_4 uFenceRegisters_28 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[28><3] , 
        \fence_regs_wr_cta_id[28><2] , \fence_regs_wr_cta_id[28><1] , 
        \fence_regs_wr_cta_id[28><0] }), .cta_id_ld(fence_regs_cta_id_ld[28]), 
        .fence_en_in(n59), .fence_en_ld(n29), .cta_id_out({
        \fence_regs_rd_cta_id[28><3] , \fence_regs_rd_cta_id[28><2] , 
        \fence_regs_rd_cta_id[28><1] , \fence_regs_rd_cta_id[28><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[28]) );
  fence_registers_1_3 uFenceRegisters_29 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[29><3] , 
        \fence_regs_wr_cta_id[29><2] , \fence_regs_wr_cta_id[29><1] , 
        \fence_regs_wr_cta_id[29><0] }), .cta_id_ld(fence_regs_cta_id_ld[29]), 
        .fence_en_in(n60), .fence_en_ld(n30), .cta_id_out({
        \fence_regs_rd_cta_id[29><3] , \fence_regs_rd_cta_id[29><2] , 
        \fence_regs_rd_cta_id[29><1] , \fence_regs_rd_cta_id[29><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[29]) );
  fence_registers_1_2 uFenceRegisters_30 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[30><3] , 
        \fence_regs_wr_cta_id[30><2] , \fence_regs_wr_cta_id[30><1] , 
        \fence_regs_wr_cta_id[30><0] }), .cta_id_ld(fence_regs_cta_id_ld[30]), 
        .fence_en_in(n64), .fence_en_ld(n31), .cta_id_out({
        \fence_regs_rd_cta_id[30><3] , \fence_regs_rd_cta_id[30><2] , 
        \fence_regs_rd_cta_id[30><1] , \fence_regs_rd_cta_id[30><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[30]) );
  fence_registers_1_1 uFenceRegisters_31 ( .clk_in(clk_in), .host_reset(n248), 
        .cta_id_in({\fence_regs_wr_cta_id[31><3] , 
        \fence_regs_wr_cta_id[31><2] , \fence_regs_wr_cta_id[31><1] , 
        \fence_regs_wr_cta_id[31><0] }), .cta_id_ld(fence_regs_cta_id_ld[31]), 
        .fence_en_in(n61), .fence_en_ld(n32), .cta_id_out({
        \fence_regs_rd_cta_id[31><3] , \fence_regs_rd_cta_id[31><2] , 
        \fence_regs_rd_cta_id[31><1] , \fence_regs_rd_cta_id[31><0] }), 
        .fence_en_out(fence_regs_rd_fence_en[31]) );
  AND2_X1 U3 ( .A1(warp_checker_fence_regs_wr_fence_en[1]), .A2(n221), .ZN(n33) );
  AND2_X1 U4 ( .A1(warp_checker_fence_regs_wr_fence_en[2]), .A2(n221), .ZN(n34) );
  AND2_X1 U5 ( .A1(warp_checker_fence_regs_wr_fence_en[4]), .A2(n222), .ZN(n35) );
  AND2_X1 U6 ( .A1(warp_checker_fence_regs_wr_fence_en[5]), .A2(n223), .ZN(n36) );
  AND2_X1 U7 ( .A1(warp_checker_fence_regs_wr_fence_en[6]), .A2(n223), .ZN(n37) );
  AND2_X1 U8 ( .A1(warp_checker_fence_regs_wr_fence_en[7]), .A2(n222), .ZN(n38) );
  AND2_X1 U9 ( .A1(warp_checker_fence_regs_wr_fence_en[8]), .A2(n222), .ZN(n39) );
  AND2_X1 U10 ( .A1(warp_checker_fence_regs_wr_fence_en[10]), .A2(n222), .ZN(
        n40) );
  AND2_X1 U11 ( .A1(warp_checker_fence_regs_wr_fence_en[11]), .A2(n222), .ZN(
        n41) );
  AND2_X1 U12 ( .A1(warp_checker_fence_regs_wr_fence_en[13]), .A2(n222), .ZN(
        n42) );
  AND2_X1 U13 ( .A1(warp_checker_fence_regs_wr_fence_en[14]), .A2(n222), .ZN(
        n43) );
  AND2_X1 U14 ( .A1(warp_checker_fence_regs_wr_fence_en[16]), .A2(n223), .ZN(
        n44) );
  AND2_X1 U15 ( .A1(warp_checker_fence_regs_wr_fence_en[18]), .A2(n225), .ZN(
        n45) );
  AND2_X1 U16 ( .A1(warp_checker_fence_regs_wr_fence_en[19]), .A2(n225), .ZN(
        n46) );
  AND2_X1 U17 ( .A1(warp_checker_fence_regs_wr_fence_en[20]), .A2(n223), .ZN(
        n47) );
  AND2_X1 U18 ( .A1(warp_checker_fence_regs_wr_fence_en[21]), .A2(n225), .ZN(
        n48) );
  AND2_X1 U19 ( .A1(warp_checker_fence_regs_wr_fence_en[22]), .A2(n225), .ZN(
        n49) );
  AND2_X1 U20 ( .A1(warp_checker_fence_regs_wr_fence_en[23]), .A2(n223), .ZN(
        n50) );
  AND2_X1 U21 ( .A1(warp_checker_fence_regs_wr_fence_en[24]), .A2(n225), .ZN(
        n51) );
  AND2_X1 U22 ( .A1(warp_checker_fence_regs_wr_fence_en[25]), .A2(n223), .ZN(
        n52) );
  AND2_X1 U23 ( .A1(warp_checker_fence_regs_wr_fence_en[26]), .A2(n225), .ZN(
        n53) );
  AND2_X1 U24 ( .A1(warp_checker_fence_regs_wr_fence_en[27]), .A2(n225), .ZN(
        n54) );
  AND2_X1 U25 ( .A1(warp_checker_fence_regs_wr_fence_en[0]), .A2(n223), .ZN(
        n55) );
  AND2_X1 U26 ( .A1(warp_checker_fence_regs_wr_fence_en[3]), .A2(n224), .ZN(
        n56) );
  AND2_X1 U27 ( .A1(warp_checker_fence_regs_wr_fence_en[9]), .A2(n224), .ZN(
        n57) );
  AND2_X1 U28 ( .A1(warp_checker_fence_regs_wr_fence_en[15]), .A2(n224), .ZN(
        n58) );
  AND2_X1 U29 ( .A1(warp_checker_fence_regs_wr_fence_en[28]), .A2(n224), .ZN(
        n59) );
  AND2_X1 U30 ( .A1(warp_checker_fence_regs_wr_fence_en[29]), .A2(n224), .ZN(
        n60) );
  AND2_X1 U31 ( .A1(warp_checker_fence_regs_wr_fence_en[31]), .A2(n224), .ZN(
        n61) );
  AND2_X1 U32 ( .A1(warp_checker_fence_regs_wr_fence_en[12]), .A2(n226), .ZN(
        n62) );
  AND2_X1 U33 ( .A1(warp_checker_fence_regs_wr_fence_en[17]), .A2(n226), .ZN(
        n63) );
  AND2_X1 U34 ( .A1(warp_checker_fence_regs_wr_fence_en[30]), .A2(n226), .ZN(
        n64) );
  INV_X1 U35 ( .A(n220), .ZN(n164) );
  INV_X1 U36 ( .A(n219), .ZN(n175) );
  INV_X1 U37 ( .A(n219), .ZN(n163) );
  INV_X1 U38 ( .A(n218), .ZN(n160) );
  INV_X1 U39 ( .A(n219), .ZN(n172) );
  INV_X1 U40 ( .A(n220), .ZN(n170) );
  INV_X1 U41 ( .A(n220), .ZN(n171) );
  INV_X1 U42 ( .A(n219), .ZN(n174) );
  INV_X1 U43 ( .A(n218), .ZN(n165) );
  INV_X1 U44 ( .A(n218), .ZN(n167) );
  INV_X1 U45 ( .A(n221), .ZN(n178) );
  INV_X1 U46 ( .A(n221), .ZN(n177) );
  BUF_X1 U47 ( .A(n229), .Z(n218) );
  BUF_X1 U48 ( .A(n237), .Z(n189) );
  BUF_X1 U49 ( .A(n232), .Z(n204) );
  BUF_X1 U50 ( .A(n235), .Z(n196) );
  BUF_X1 U51 ( .A(n234), .Z(n197) );
  BUF_X1 U52 ( .A(n237), .Z(n190) );
  BUF_X1 U53 ( .A(n235), .Z(n194) );
  BUF_X1 U54 ( .A(n236), .Z(n193) );
  BUF_X1 U55 ( .A(n236), .Z(n192) );
  BUF_X1 U56 ( .A(n230), .Z(n210) );
  BUF_X1 U57 ( .A(n230), .Z(n217) );
  BUF_X1 U58 ( .A(n230), .Z(n216) );
  BUF_X1 U59 ( .A(n235), .Z(n195) );
  BUF_X1 U60 ( .A(n236), .Z(n191) );
  BUF_X1 U61 ( .A(n231), .Z(n209) );
  BUF_X1 U62 ( .A(n234), .Z(n199) );
  BUF_X1 U63 ( .A(n234), .Z(n198) );
  BUF_X1 U64 ( .A(n231), .Z(n207) );
  BUF_X1 U65 ( .A(n231), .Z(n206) );
  BUF_X1 U66 ( .A(n232), .Z(n205) );
  BUF_X1 U67 ( .A(n233), .Z(n202) );
  BUF_X1 U68 ( .A(n233), .Z(n201) );
  BUF_X1 U69 ( .A(n233), .Z(n200) );
  BUF_X1 U70 ( .A(n232), .Z(n203) );
  BUF_X1 U71 ( .A(n229), .Z(n220) );
  BUF_X1 U72 ( .A(n229), .Z(n219) );
  BUF_X1 U73 ( .A(n228), .Z(n221) );
  BUF_X1 U74 ( .A(n238), .Z(n186) );
  BUF_X1 U75 ( .A(n239), .Z(n183) );
  BUF_X1 U76 ( .A(n238), .Z(n187) );
  BUF_X1 U77 ( .A(n239), .Z(n182) );
  BUF_X1 U78 ( .A(n239), .Z(n184) );
  BUF_X1 U79 ( .A(n237), .Z(n188) );
  BUF_X1 U80 ( .A(n238), .Z(n185) );
  BUF_X1 U81 ( .A(n240), .Z(n181) );
  BUF_X1 U82 ( .A(n228), .Z(n222) );
  BUF_X1 U83 ( .A(n227), .Z(n225) );
  BUF_X1 U84 ( .A(n227), .Z(n224) );
  BUF_X1 U85 ( .A(n228), .Z(n223) );
  BUF_X1 U86 ( .A(n227), .Z(n226) );
  BUF_X1 U87 ( .A(n240), .Z(n179) );
  BUF_X1 U88 ( .A(n240), .Z(n180) );
  BUF_X1 U89 ( .A(n244), .Z(n234) );
  BUF_X1 U90 ( .A(n243), .Z(n235) );
  BUF_X1 U91 ( .A(n243), .Z(n236) );
  BUF_X1 U92 ( .A(n242), .Z(n237) );
  BUF_X1 U93 ( .A(n244), .Z(n233) );
  BUF_X1 U94 ( .A(n246), .Z(n230) );
  BUF_X1 U95 ( .A(n245), .Z(n231) );
  BUF_X1 U96 ( .A(n245), .Z(n232) );
  BUF_X1 U97 ( .A(n246), .Z(n229) );
  BUF_X1 U98 ( .A(n241), .Z(n239) );
  BUF_X1 U99 ( .A(n242), .Z(n238) );
  BUF_X1 U100 ( .A(n241), .Z(n240) );
  BUF_X1 U101 ( .A(n247), .Z(n227) );
  BUF_X1 U102 ( .A(n247), .Z(n228) );
  INV_X1 U103 ( .A(n158), .ZN(n244) );
  INV_X1 U104 ( .A(n158), .ZN(n243) );
  INV_X1 U105 ( .A(n158), .ZN(n242) );
  INV_X1 U106 ( .A(n159), .ZN(n246) );
  INV_X1 U107 ( .A(n159), .ZN(n245) );
  INV_X1 U108 ( .A(n158), .ZN(n241) );
  INV_X1 U109 ( .A(n159), .ZN(n247) );
  BUF_X1 U110 ( .A(warp_scheduler_reset), .Z(n158) );
  BUF_X1 U111 ( .A(warp_scheduler_reset), .Z(n159) );
  AND2_X1 U112 ( .A1(fence_regs_rd_fence_en[1]), .A2(n201), .ZN(
        warp_checker_fence_regs_rd_fence_en[1]) );
  AND2_X1 U113 ( .A1(fence_regs_rd_fence_en[0]), .A2(n199), .ZN(
        warp_checker_fence_regs_rd_fence_en[0]) );
  AND2_X1 U114 ( .A1(fence_regs_rd_fence_en[22]), .A2(n201), .ZN(
        warp_checker_fence_regs_rd_fence_en[22]) );
  AND2_X1 U115 ( .A1(fence_regs_rd_fence_en[18]), .A2(n201), .ZN(
        warp_checker_fence_regs_rd_fence_en[18]) );
  AND2_X1 U116 ( .A1(fence_regs_rd_fence_en[14]), .A2(n200), .ZN(
        warp_checker_fence_regs_rd_fence_en[14]) );
  AND2_X1 U117 ( .A1(fence_regs_rd_fence_en[9]), .A2(n189), .ZN(
        warp_checker_fence_regs_rd_fence_en[9]) );
  AND2_X1 U118 ( .A1(fence_regs_rd_fence_en[26]), .A2(n202), .ZN(
        warp_checker_fence_regs_rd_fence_en[26]) );
  AND2_X1 U119 ( .A1(fence_regs_rd_fence_en[30]), .A2(n203), .ZN(
        warp_checker_fence_regs_rd_fence_en[30]) );
  AND2_X1 U120 ( .A1(fence_regs_rd_fence_en[31]), .A2(n203), .ZN(
        warp_checker_fence_regs_rd_fence_en[31]) );
  AND2_X1 U121 ( .A1(fence_regs_rd_fence_en[2]), .A2(n203), .ZN(
        warp_checker_fence_regs_rd_fence_en[2]) );
  AND2_X1 U122 ( .A1(fence_regs_rd_fence_en[16]), .A2(n200), .ZN(
        warp_checker_fence_regs_rd_fence_en[16]) );
  AND2_X1 U123 ( .A1(fence_regs_rd_fence_en[15]), .A2(n200), .ZN(
        warp_checker_fence_regs_rd_fence_en[15]) );
  AND2_X1 U124 ( .A1(fence_regs_rd_fence_en[11]), .A2(n200), .ZN(
        warp_checker_fence_regs_rd_fence_en[11]) );
  AND2_X1 U125 ( .A1(fence_regs_rd_fence_en[23]), .A2(n202), .ZN(
        warp_checker_fence_regs_rd_fence_en[23]) );
  AND2_X1 U126 ( .A1(fence_regs_rd_fence_en[19]), .A2(n201), .ZN(
        warp_checker_fence_regs_rd_fence_en[19]) );
  AND2_X1 U127 ( .A1(fence_regs_rd_fence_en[29]), .A2(n202), .ZN(
        warp_checker_fence_regs_rd_fence_en[29]) );
  AND2_X1 U128 ( .A1(fence_regs_rd_fence_en[28]), .A2(n202), .ZN(
        warp_checker_fence_regs_rd_fence_en[28]) );
  AND2_X1 U129 ( .A1(fence_regs_rd_fence_en[27]), .A2(n202), .ZN(
        warp_checker_fence_regs_rd_fence_en[27]) );
  AND2_X1 U130 ( .A1(fence_regs_rd_fence_en[17]), .A2(n201), .ZN(
        warp_checker_fence_regs_rd_fence_en[17]) );
  AND2_X1 U131 ( .A1(fence_regs_rd_fence_en[7]), .A2(n204), .ZN(
        warp_checker_fence_regs_rd_fence_en[7]) );
  AND2_X1 U132 ( .A1(fence_regs_rd_fence_en[10]), .A2(n200), .ZN(
        warp_checker_fence_regs_rd_fence_en[10]) );
  AND2_X1 U133 ( .A1(fence_regs_rd_fence_en[13]), .A2(n200), .ZN(
        warp_checker_fence_regs_rd_fence_en[13]) );
  AND2_X1 U134 ( .A1(fence_regs_rd_fence_en[12]), .A2(n200), .ZN(
        warp_checker_fence_regs_rd_fence_en[12]) );
  AND2_X1 U135 ( .A1(fence_regs_rd_fence_en[25]), .A2(n202), .ZN(
        warp_checker_fence_regs_rd_fence_en[25]) );
  AND2_X1 U136 ( .A1(fence_regs_rd_fence_en[24]), .A2(n202), .ZN(
        warp_checker_fence_regs_rd_fence_en[24]) );
  AND2_X1 U137 ( .A1(fence_regs_rd_fence_en[21]), .A2(n201), .ZN(
        warp_checker_fence_regs_rd_fence_en[21]) );
  AND2_X1 U138 ( .A1(fence_regs_rd_fence_en[20]), .A2(n201), .ZN(
        warp_checker_fence_regs_rd_fence_en[20]) );
  AND2_X1 U139 ( .A1(fence_regs_rd_fence_en[8]), .A2(n204), .ZN(
        warp_checker_fence_regs_rd_fence_en[8]) );
  AND2_X1 U140 ( .A1(fence_regs_rd_fence_en[3]), .A2(n203), .ZN(
        warp_checker_fence_regs_rd_fence_en[3]) );
  AND2_X1 U141 ( .A1(fence_regs_rd_fence_en[4]), .A2(n203), .ZN(
        warp_checker_fence_regs_rd_fence_en[4]) );
  AND2_X1 U142 ( .A1(\fence_regs_rd_cta_id[21><2] ), .A2(n218), .ZN(
        \warp_checker_fence_regs_rd_cta_id[21><2] ) );
  AND2_X1 U143 ( .A1(fence_regs_rd_fence_en[5]), .A2(n203), .ZN(
        warp_checker_fence_regs_rd_fence_en[5]) );
  AND2_X1 U144 ( .A1(fence_regs_rd_fence_en[6]), .A2(n203), .ZN(
        warp_checker_fence_regs_rd_fence_en[6]) );
  AND2_X1 U145 ( .A1(\fence_regs_rd_cta_id[22><1] ), .A2(n218), .ZN(
        \warp_checker_fence_regs_rd_cta_id[22><1] ) );
  AND2_X1 U146 ( .A1(\fence_regs_rd_cta_id[22><0] ), .A2(n218), .ZN(
        \warp_checker_fence_regs_rd_cta_id[22><0] ) );
  AND2_X1 U147 ( .A1(\fence_regs_rd_cta_id[21><3] ), .A2(n218), .ZN(
        \warp_checker_fence_regs_rd_cta_id[21><3] ) );
  AND2_X1 U148 ( .A1(\fence_regs_rd_cta_id[23><1] ), .A2(n189), .ZN(
        \warp_checker_fence_regs_rd_cta_id[23><1] ) );
  AND2_X1 U149 ( .A1(\fence_regs_rd_cta_id[0><1] ), .A2(n204), .ZN(
        \warp_checker_fence_regs_rd_cta_id[0><1] ) );
  AND2_X1 U150 ( .A1(\fence_regs_rd_cta_id[0><2] ), .A2(n204), .ZN(
        \warp_checker_fence_regs_rd_cta_id[0><2] ) );
  AND2_X1 U151 ( .A1(\fence_regs_rd_cta_id[0><3] ), .A2(n204), .ZN(
        \warp_checker_fence_regs_rd_cta_id[0><3] ) );
  AND2_X1 U152 ( .A1(\fence_regs_rd_cta_id[5><1] ), .A2(n197), .ZN(
        \warp_checker_fence_regs_rd_cta_id[5><1] ) );
  AND2_X1 U153 ( .A1(\fence_regs_rd_cta_id[5><2] ), .A2(n197), .ZN(
        \warp_checker_fence_regs_rd_cta_id[5><2] ) );
  AND2_X1 U154 ( .A1(\fence_regs_rd_cta_id[5><3] ), .A2(n197), .ZN(
        \warp_checker_fence_regs_rd_cta_id[5><3] ) );
  AND2_X1 U155 ( .A1(\fence_regs_rd_cta_id[4><1] ), .A2(n196), .ZN(
        \warp_checker_fence_regs_rd_cta_id[4><1] ) );
  AND2_X1 U156 ( .A1(\fence_regs_rd_cta_id[4><2] ), .A2(n196), .ZN(
        \warp_checker_fence_regs_rd_cta_id[4><2] ) );
  AND2_X1 U157 ( .A1(\fence_regs_rd_cta_id[4><3] ), .A2(n196), .ZN(
        \warp_checker_fence_regs_rd_cta_id[4><3] ) );
  AND2_X1 U158 ( .A1(\fence_regs_rd_cta_id[9><1] ), .A2(n199), .ZN(
        \warp_checker_fence_regs_rd_cta_id[9><1] ) );
  AND2_X1 U159 ( .A1(\fence_regs_rd_cta_id[9><2] ), .A2(n199), .ZN(
        \warp_checker_fence_regs_rd_cta_id[9><2] ) );
  AND2_X1 U160 ( .A1(\fence_regs_rd_cta_id[9><3] ), .A2(n199), .ZN(
        \warp_checker_fence_regs_rd_cta_id[9><3] ) );
  AND2_X1 U161 ( .A1(\fence_regs_rd_cta_id[0><0] ), .A2(n204), .ZN(
        \warp_checker_fence_regs_rd_cta_id[0><0] ) );
  AND2_X1 U162 ( .A1(\fence_regs_rd_cta_id[5><0] ), .A2(n197), .ZN(
        \warp_checker_fence_regs_rd_cta_id[5><0] ) );
  AND2_X1 U163 ( .A1(\fence_regs_rd_cta_id[4><0] ), .A2(n196), .ZN(
        \warp_checker_fence_regs_rd_cta_id[4><0] ) );
  AND2_X1 U164 ( .A1(\fence_regs_rd_cta_id[9><0] ), .A2(n199), .ZN(
        \warp_checker_fence_regs_rd_cta_id[9><0] ) );
  AND2_X1 U165 ( .A1(\fence_regs_rd_cta_id[3><1] ), .A2(n193), .ZN(
        \warp_checker_fence_regs_rd_cta_id[3><1] ) );
  AND2_X1 U166 ( .A1(\fence_regs_rd_cta_id[3><2] ), .A2(n196), .ZN(
        \warp_checker_fence_regs_rd_cta_id[3><2] ) );
  AND2_X1 U167 ( .A1(\fence_regs_rd_cta_id[3><3] ), .A2(n196), .ZN(
        \warp_checker_fence_regs_rd_cta_id[3><3] ) );
  AND2_X1 U168 ( .A1(\fence_regs_rd_cta_id[6><1] ), .A2(n197), .ZN(
        \warp_checker_fence_regs_rd_cta_id[6><1] ) );
  AND2_X1 U169 ( .A1(\fence_regs_rd_cta_id[6><2] ), .A2(n197), .ZN(
        \warp_checker_fence_regs_rd_cta_id[6><2] ) );
  AND2_X1 U170 ( .A1(\fence_regs_rd_cta_id[6><3] ), .A2(n198), .ZN(
        \warp_checker_fence_regs_rd_cta_id[6><3] ) );
  AND2_X1 U171 ( .A1(\fence_regs_rd_cta_id[14><1] ), .A2(n207), .ZN(
        \warp_checker_fence_regs_rd_cta_id[14><1] ) );
  AND2_X1 U172 ( .A1(\fence_regs_rd_cta_id[14><2] ), .A2(n207), .ZN(
        \warp_checker_fence_regs_rd_cta_id[14><2] ) );
  AND2_X1 U173 ( .A1(\fence_regs_rd_cta_id[14><3] ), .A2(n207), .ZN(
        \warp_checker_fence_regs_rd_cta_id[14><3] ) );
  AND2_X1 U174 ( .A1(\fence_regs_rd_cta_id[26><1] ), .A2(n191), .ZN(
        \warp_checker_fence_regs_rd_cta_id[26><1] ) );
  AND2_X1 U175 ( .A1(\fence_regs_rd_cta_id[26><2] ), .A2(n191), .ZN(
        \warp_checker_fence_regs_rd_cta_id[26><2] ) );
  AND2_X1 U176 ( .A1(\fence_regs_rd_cta_id[26><3] ), .A2(n194), .ZN(
        \warp_checker_fence_regs_rd_cta_id[26><3] ) );
  AND2_X1 U177 ( .A1(\fence_regs_rd_cta_id[30><1] ), .A2(n192), .ZN(
        \warp_checker_fence_regs_rd_cta_id[30><1] ) );
  AND2_X1 U178 ( .A1(\fence_regs_rd_cta_id[30><2] ), .A2(n194), .ZN(
        \warp_checker_fence_regs_rd_cta_id[30><2] ) );
  AND2_X1 U179 ( .A1(\fence_regs_rd_cta_id[30><3] ), .A2(n193), .ZN(
        \warp_checker_fence_regs_rd_cta_id[30><3] ) );
  AND2_X1 U180 ( .A1(\fence_regs_rd_cta_id[22><2] ), .A2(n196), .ZN(
        \warp_checker_fence_regs_rd_cta_id[22><2] ) );
  AND2_X1 U181 ( .A1(\fence_regs_rd_cta_id[22><3] ), .A2(n192), .ZN(
        \warp_checker_fence_regs_rd_cta_id[22><3] ) );
  AND2_X1 U182 ( .A1(\fence_regs_rd_cta_id[18><1] ), .A2(n210), .ZN(
        \warp_checker_fence_regs_rd_cta_id[18><1] ) );
  AND2_X1 U183 ( .A1(\fence_regs_rd_cta_id[18><2] ), .A2(n210), .ZN(
        \warp_checker_fence_regs_rd_cta_id[18><2] ) );
  AND2_X1 U184 ( .A1(\fence_regs_rd_cta_id[18><3] ), .A2(n216), .ZN(
        \warp_checker_fence_regs_rd_cta_id[18><3] ) );
  AND2_X1 U185 ( .A1(\fence_regs_rd_cta_id[3><0] ), .A2(n195), .ZN(
        \warp_checker_fence_regs_rd_cta_id[3><0] ) );
  AND2_X1 U186 ( .A1(\fence_regs_rd_cta_id[6><0] ), .A2(n197), .ZN(
        \warp_checker_fence_regs_rd_cta_id[6><0] ) );
  AND2_X1 U187 ( .A1(\fence_regs_rd_cta_id[14><0] ), .A2(n207), .ZN(
        \warp_checker_fence_regs_rd_cta_id[14><0] ) );
  AND2_X1 U188 ( .A1(\fence_regs_rd_cta_id[26><0] ), .A2(n190), .ZN(
        \warp_checker_fence_regs_rd_cta_id[26><0] ) );
  AND2_X1 U189 ( .A1(\fence_regs_rd_cta_id[30><0] ), .A2(n192), .ZN(
        \warp_checker_fence_regs_rd_cta_id[30><0] ) );
  AND2_X1 U190 ( .A1(\fence_regs_rd_cta_id[18><0] ), .A2(n210), .ZN(
        \warp_checker_fence_regs_rd_cta_id[18><0] ) );
  AND2_X1 U191 ( .A1(\fence_regs_rd_cta_id[1><1] ), .A2(n216), .ZN(
        \warp_checker_fence_regs_rd_cta_id[1><1] ) );
  AND2_X1 U192 ( .A1(\fence_regs_rd_cta_id[1><2] ), .A2(n216), .ZN(
        \warp_checker_fence_regs_rd_cta_id[1><2] ) );
  AND2_X1 U193 ( .A1(\fence_regs_rd_cta_id[1><3] ), .A2(n217), .ZN(
        \warp_checker_fence_regs_rd_cta_id[1><3] ) );
  AND2_X1 U194 ( .A1(\fence_regs_rd_cta_id[25><1] ), .A2(n190), .ZN(
        \warp_checker_fence_regs_rd_cta_id[25><1] ) );
  AND2_X1 U195 ( .A1(\fence_regs_rd_cta_id[25><2] ), .A2(n190), .ZN(
        \warp_checker_fence_regs_rd_cta_id[25><2] ) );
  AND2_X1 U196 ( .A1(\fence_regs_rd_cta_id[25><3] ), .A2(n194), .ZN(
        \warp_checker_fence_regs_rd_cta_id[25><3] ) );
  AND2_X1 U197 ( .A1(\fence_regs_rd_cta_id[24><1] ), .A2(n193), .ZN(
        \warp_checker_fence_regs_rd_cta_id[24><1] ) );
  AND2_X1 U198 ( .A1(\fence_regs_rd_cta_id[24><2] ), .A2(n190), .ZN(
        \warp_checker_fence_regs_rd_cta_id[24><2] ) );
  AND2_X1 U199 ( .A1(\fence_regs_rd_cta_id[24><3] ), .A2(n190), .ZN(
        \warp_checker_fence_regs_rd_cta_id[24><3] ) );
  AND2_X1 U200 ( .A1(\fence_regs_rd_cta_id[23><2] ), .A2(n193), .ZN(
        \warp_checker_fence_regs_rd_cta_id[23><2] ) );
  AND2_X1 U201 ( .A1(\fence_regs_rd_cta_id[23><3] ), .A2(n190), .ZN(
        \warp_checker_fence_regs_rd_cta_id[23><3] ) );
  AND2_X1 U202 ( .A1(\fence_regs_rd_cta_id[21><0] ), .A2(n217), .ZN(
        \warp_checker_fence_regs_rd_cta_id[21><0] ) );
  AND2_X1 U203 ( .A1(\fence_regs_rd_cta_id[21><1] ), .A2(n217), .ZN(
        \warp_checker_fence_regs_rd_cta_id[21><1] ) );
  AND2_X1 U204 ( .A1(\fence_regs_rd_cta_id[20><1] ), .A2(n217), .ZN(
        \warp_checker_fence_regs_rd_cta_id[20><1] ) );
  AND2_X1 U205 ( .A1(\fence_regs_rd_cta_id[20><2] ), .A2(n217), .ZN(
        \warp_checker_fence_regs_rd_cta_id[20><2] ) );
  AND2_X1 U206 ( .A1(\fence_regs_rd_cta_id[20><3] ), .A2(n217), .ZN(
        \warp_checker_fence_regs_rd_cta_id[20><3] ) );
  AND2_X1 U207 ( .A1(\fence_regs_rd_cta_id[19><1] ), .A2(n209), .ZN(
        \warp_checker_fence_regs_rd_cta_id[19><1] ) );
  AND2_X1 U208 ( .A1(\fence_regs_rd_cta_id[19><2] ), .A2(n216), .ZN(
        \warp_checker_fence_regs_rd_cta_id[19><2] ) );
  AND2_X1 U209 ( .A1(\fence_regs_rd_cta_id[19><3] ), .A2(n216), .ZN(
        \warp_checker_fence_regs_rd_cta_id[19><3] ) );
  AND2_X1 U210 ( .A1(\fence_regs_rd_cta_id[29><1] ), .A2(n195), .ZN(
        \warp_checker_fence_regs_rd_cta_id[29><1] ) );
  AND2_X1 U211 ( .A1(\fence_regs_rd_cta_id[29><2] ), .A2(n192), .ZN(
        \warp_checker_fence_regs_rd_cta_id[29><2] ) );
  AND2_X1 U212 ( .A1(\fence_regs_rd_cta_id[29><3] ), .A2(n192), .ZN(
        \warp_checker_fence_regs_rd_cta_id[29><3] ) );
  AND2_X1 U213 ( .A1(\fence_regs_rd_cta_id[28><1] ), .A2(n191), .ZN(
        \warp_checker_fence_regs_rd_cta_id[28><1] ) );
  AND2_X1 U214 ( .A1(\fence_regs_rd_cta_id[28><2] ), .A2(n194), .ZN(
        \warp_checker_fence_regs_rd_cta_id[28><2] ) );
  AND2_X1 U215 ( .A1(\fence_regs_rd_cta_id[28><3] ), .A2(n195), .ZN(
        \warp_checker_fence_regs_rd_cta_id[28><3] ) );
  AND2_X1 U216 ( .A1(\fence_regs_rd_cta_id[27><1] ), .A2(n191), .ZN(
        \warp_checker_fence_regs_rd_cta_id[27><1] ) );
  AND2_X1 U217 ( .A1(\fence_regs_rd_cta_id[27><2] ), .A2(n191), .ZN(
        \warp_checker_fence_regs_rd_cta_id[27><2] ) );
  AND2_X1 U218 ( .A1(\fence_regs_rd_cta_id[27><3] ), .A2(n194), .ZN(
        \warp_checker_fence_regs_rd_cta_id[27><3] ) );
  AND2_X1 U219 ( .A1(\fence_regs_rd_cta_id[17><1] ), .A2(n210), .ZN(
        \warp_checker_fence_regs_rd_cta_id[17><1] ) );
  AND2_X1 U220 ( .A1(\fence_regs_rd_cta_id[17><2] ), .A2(n210), .ZN(
        \warp_checker_fence_regs_rd_cta_id[17><2] ) );
  AND2_X1 U221 ( .A1(\fence_regs_rd_cta_id[17><3] ), .A2(n210), .ZN(
        \warp_checker_fence_regs_rd_cta_id[17><3] ) );
  AND2_X1 U222 ( .A1(\fence_regs_rd_cta_id[16><1] ), .A2(n209), .ZN(
        \warp_checker_fence_regs_rd_cta_id[16><1] ) );
  AND2_X1 U223 ( .A1(\fence_regs_rd_cta_id[16><2] ), .A2(n209), .ZN(
        \warp_checker_fence_regs_rd_cta_id[16><2] ) );
  AND2_X1 U224 ( .A1(\fence_regs_rd_cta_id[16><3] ), .A2(n209), .ZN(
        \warp_checker_fence_regs_rd_cta_id[16><3] ) );
  AND2_X1 U225 ( .A1(\fence_regs_rd_cta_id[15><1] ), .A2(n207), .ZN(
        \warp_checker_fence_regs_rd_cta_id[15><1] ) );
  AND2_X1 U226 ( .A1(\fence_regs_rd_cta_id[15><2] ), .A2(n209), .ZN(
        \warp_checker_fence_regs_rd_cta_id[15><2] ) );
  AND2_X1 U227 ( .A1(\fence_regs_rd_cta_id[15><3] ), .A2(n209), .ZN(
        \warp_checker_fence_regs_rd_cta_id[15><3] ) );
  AND2_X1 U228 ( .A1(\fence_regs_rd_cta_id[10><1] ), .A2(n205), .ZN(
        \warp_checker_fence_regs_rd_cta_id[10><1] ) );
  AND2_X1 U229 ( .A1(\fence_regs_rd_cta_id[10><2] ), .A2(n205), .ZN(
        \warp_checker_fence_regs_rd_cta_id[10><2] ) );
  AND2_X1 U230 ( .A1(\fence_regs_rd_cta_id[10><3] ), .A2(n205), .ZN(
        \warp_checker_fence_regs_rd_cta_id[10><3] ) );
  AND2_X1 U231 ( .A1(\fence_regs_rd_cta_id[8><1] ), .A2(n198), .ZN(
        \warp_checker_fence_regs_rd_cta_id[8><1] ) );
  AND2_X1 U232 ( .A1(\fence_regs_rd_cta_id[8><2] ), .A2(n199), .ZN(
        \warp_checker_fence_regs_rd_cta_id[8><2] ) );
  AND2_X1 U233 ( .A1(\fence_regs_rd_cta_id[8><3] ), .A2(n199), .ZN(
        \warp_checker_fence_regs_rd_cta_id[8><3] ) );
  AND2_X1 U234 ( .A1(\fence_regs_rd_cta_id[7><1] ), .A2(n198), .ZN(
        \warp_checker_fence_regs_rd_cta_id[7><1] ) );
  AND2_X1 U235 ( .A1(\fence_regs_rd_cta_id[7><2] ), .A2(n198), .ZN(
        \warp_checker_fence_regs_rd_cta_id[7><2] ) );
  AND2_X1 U236 ( .A1(\fence_regs_rd_cta_id[7><3] ), .A2(n198), .ZN(
        \warp_checker_fence_regs_rd_cta_id[7><3] ) );
  AND2_X1 U237 ( .A1(\fence_regs_rd_cta_id[13><1] ), .A2(n206), .ZN(
        \warp_checker_fence_regs_rd_cta_id[13><1] ) );
  AND2_X1 U238 ( .A1(\fence_regs_rd_cta_id[13><2] ), .A2(n206), .ZN(
        \warp_checker_fence_regs_rd_cta_id[13><2] ) );
  AND2_X1 U239 ( .A1(\fence_regs_rd_cta_id[13><3] ), .A2(n207), .ZN(
        \warp_checker_fence_regs_rd_cta_id[13><3] ) );
  AND2_X1 U240 ( .A1(\fence_regs_rd_cta_id[12><1] ), .A2(n206), .ZN(
        \warp_checker_fence_regs_rd_cta_id[12><1] ) );
  AND2_X1 U241 ( .A1(\fence_regs_rd_cta_id[12><2] ), .A2(n206), .ZN(
        \warp_checker_fence_regs_rd_cta_id[12><2] ) );
  AND2_X1 U242 ( .A1(\fence_regs_rd_cta_id[12><3] ), .A2(n206), .ZN(
        \warp_checker_fence_regs_rd_cta_id[12><3] ) );
  AND2_X1 U243 ( .A1(\fence_regs_rd_cta_id[11><1] ), .A2(n205), .ZN(
        \warp_checker_fence_regs_rd_cta_id[11><1] ) );
  AND2_X1 U244 ( .A1(\fence_regs_rd_cta_id[11><2] ), .A2(n205), .ZN(
        \warp_checker_fence_regs_rd_cta_id[11><2] ) );
  AND2_X1 U245 ( .A1(\fence_regs_rd_cta_id[11><3] ), .A2(n205), .ZN(
        \warp_checker_fence_regs_rd_cta_id[11><3] ) );
  AND2_X1 U246 ( .A1(\fence_regs_rd_cta_id[1><0] ), .A2(n216), .ZN(
        \warp_checker_fence_regs_rd_cta_id[1><0] ) );
  AND2_X1 U247 ( .A1(\fence_regs_rd_cta_id[2><1] ), .A2(n192), .ZN(
        \warp_checker_fence_regs_rd_cta_id[2><1] ) );
  AND2_X1 U248 ( .A1(\fence_regs_rd_cta_id[2><2] ), .A2(n192), .ZN(
        \warp_checker_fence_regs_rd_cta_id[2><2] ) );
  AND2_X1 U249 ( .A1(\fence_regs_rd_cta_id[2><3] ), .A2(n195), .ZN(
        \warp_checker_fence_regs_rd_cta_id[2><3] ) );
  AND2_X1 U250 ( .A1(\fence_regs_rd_cta_id[31><1] ), .A2(n195), .ZN(
        \warp_checker_fence_regs_rd_cta_id[31><1] ) );
  AND2_X1 U251 ( .A1(\fence_regs_rd_cta_id[31><2] ), .A2(n193), .ZN(
        \warp_checker_fence_regs_rd_cta_id[31><2] ) );
  AND2_X1 U252 ( .A1(\fence_regs_rd_cta_id[31><3] ), .A2(n195), .ZN(
        \warp_checker_fence_regs_rd_cta_id[31><3] ) );
  AND2_X1 U253 ( .A1(\fence_regs_rd_cta_id[25><0] ), .A2(n195), .ZN(
        \warp_checker_fence_regs_rd_cta_id[25><0] ) );
  AND2_X1 U254 ( .A1(\fence_regs_rd_cta_id[24><0] ), .A2(n190), .ZN(
        \warp_checker_fence_regs_rd_cta_id[24><0] ) );
  AND2_X1 U255 ( .A1(\fence_regs_rd_cta_id[23><0] ), .A2(n193), .ZN(
        \warp_checker_fence_regs_rd_cta_id[23><0] ) );
  AND2_X1 U256 ( .A1(\fence_regs_rd_cta_id[20><0] ), .A2(n217), .ZN(
        \warp_checker_fence_regs_rd_cta_id[20><0] ) );
  AND2_X1 U257 ( .A1(\fence_regs_rd_cta_id[19><0] ), .A2(n216), .ZN(
        \warp_checker_fence_regs_rd_cta_id[19><0] ) );
  AND2_X1 U258 ( .A1(\fence_regs_rd_cta_id[29><0] ), .A2(n191), .ZN(
        \warp_checker_fence_regs_rd_cta_id[29><0] ) );
  AND2_X1 U259 ( .A1(\fence_regs_rd_cta_id[28><0] ), .A2(n191), .ZN(
        \warp_checker_fence_regs_rd_cta_id[28><0] ) );
  AND2_X1 U260 ( .A1(\fence_regs_rd_cta_id[27><0] ), .A2(n194), .ZN(
        \warp_checker_fence_regs_rd_cta_id[27><0] ) );
  AND2_X1 U261 ( .A1(\fence_regs_rd_cta_id[17><0] ), .A2(n210), .ZN(
        \warp_checker_fence_regs_rd_cta_id[17><0] ) );
  AND2_X1 U262 ( .A1(\fence_regs_rd_cta_id[16><0] ), .A2(n209), .ZN(
        \warp_checker_fence_regs_rd_cta_id[16><0] ) );
  AND2_X1 U263 ( .A1(\fence_regs_rd_cta_id[15><0] ), .A2(n207), .ZN(
        \warp_checker_fence_regs_rd_cta_id[15><0] ) );
  AND2_X1 U264 ( .A1(\fence_regs_rd_cta_id[10><0] ), .A2(n204), .ZN(
        \warp_checker_fence_regs_rd_cta_id[10><0] ) );
  AND2_X1 U265 ( .A1(\fence_regs_rd_cta_id[8><0] ), .A2(n198), .ZN(
        \warp_checker_fence_regs_rd_cta_id[8><0] ) );
  AND2_X1 U266 ( .A1(\fence_regs_rd_cta_id[7><0] ), .A2(n198), .ZN(
        \warp_checker_fence_regs_rd_cta_id[7><0] ) );
  AND2_X1 U267 ( .A1(\fence_regs_rd_cta_id[13><0] ), .A2(n206), .ZN(
        \warp_checker_fence_regs_rd_cta_id[13><0] ) );
  AND2_X1 U268 ( .A1(\fence_regs_rd_cta_id[12><0] ), .A2(n206), .ZN(
        \warp_checker_fence_regs_rd_cta_id[12><0] ) );
  AND2_X1 U269 ( .A1(\fence_regs_rd_cta_id[11><0] ), .A2(n205), .ZN(
        \warp_checker_fence_regs_rd_cta_id[11><0] ) );
  AND2_X1 U270 ( .A1(\fence_regs_rd_cta_id[2><0] ), .A2(n194), .ZN(
        \warp_checker_fence_regs_rd_cta_id[2><0] ) );
  AND2_X1 U271 ( .A1(\fence_regs_rd_cta_id[31><0] ), .A2(n193), .ZN(
        \warp_checker_fence_regs_rd_cta_id[31><0] ) );
  AND2_X1 U272 ( .A1(warp_gen_fence_regs_cta_id_ld[3]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[3]) );
  AND2_X1 U273 ( .A1(warp_gen_fence_regs_cta_id_ld[4]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[4]) );
  AND2_X1 U274 ( .A1(warp_gen_fence_regs_cta_id_ld[5]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[5]) );
  AND2_X1 U275 ( .A1(warp_gen_fence_regs_cta_id_ld[6]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[6]) );
  AND2_X1 U276 ( .A1(warp_gen_fence_regs_cta_id_ld[7]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[7]) );
  AND2_X1 U277 ( .A1(warp_gen_fence_regs_cta_id_ld[8]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[8]) );
  AND2_X1 U278 ( .A1(warp_gen_fence_regs_cta_id_ld[9]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[9]) );
  AND2_X1 U279 ( .A1(warp_gen_fence_regs_cta_id_ld[30]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[30]) );
  AND2_X1 U280 ( .A1(warp_gen_fence_regs_cta_id_ld[31]), .A2(n173), .ZN(
        fence_regs_cta_id_ld[31]) );
  AND2_X1 U281 ( .A1(warp_gen_fence_regs_cta_id_ld[10]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[10]) );
  AND2_X1 U282 ( .A1(warp_gen_fence_regs_cta_id_ld[11]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[11]) );
  AND2_X1 U283 ( .A1(warp_gen_fence_regs_cta_id_ld[12]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[12]) );
  AND2_X1 U284 ( .A1(warp_gen_fence_regs_cta_id_ld[13]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[13]) );
  AND2_X1 U285 ( .A1(warp_gen_fence_regs_cta_id_ld[14]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[14]) );
  AND2_X1 U286 ( .A1(warp_gen_fence_regs_cta_id_ld[15]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[15]) );
  AND2_X1 U287 ( .A1(warp_gen_fence_regs_cta_id_ld[16]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[16]) );
  AND2_X1 U288 ( .A1(warp_gen_fence_regs_cta_id_ld[0]), .A2(n175), .ZN(
        fence_regs_cta_id_ld[0]) );
  AND2_X1 U289 ( .A1(warp_gen_fence_regs_cta_id_ld[1]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[1]) );
  AND2_X1 U290 ( .A1(warp_gen_fence_regs_cta_id_ld[2]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[2]) );
  AND2_X1 U291 ( .A1(warp_gen_fence_regs_cta_id_ld[17]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[17]) );
  AND2_X1 U292 ( .A1(warp_gen_fence_regs_cta_id_ld[18]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[18]) );
  AND2_X1 U293 ( .A1(warp_gen_fence_regs_cta_id_ld[19]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[19]) );
  AND2_X1 U294 ( .A1(warp_gen_fence_regs_cta_id_ld[20]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[20]) );
  AND2_X1 U295 ( .A1(warp_gen_fence_regs_cta_id_ld[21]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[21]) );
  AND2_X1 U296 ( .A1(warp_gen_fence_regs_cta_id_ld[22]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[22]) );
  AND2_X1 U297 ( .A1(warp_gen_fence_regs_cta_id_ld[23]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[23]) );
  AND2_X1 U298 ( .A1(warp_gen_fence_regs_cta_id_ld[24]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[24]) );
  AND2_X1 U299 ( .A1(warp_gen_fence_regs_cta_id_ld[25]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[25]) );
  AND2_X1 U300 ( .A1(warp_gen_fence_regs_cta_id_ld[26]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[26]) );
  AND2_X1 U301 ( .A1(warp_gen_fence_regs_cta_id_ld[27]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[27]) );
  AND2_X1 U302 ( .A1(warp_gen_fence_regs_cta_id_ld[28]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[28]) );
  AND2_X1 U303 ( .A1(warp_gen_fence_regs_cta_id_ld[29]), .A2(n174), .ZN(
        fence_regs_cta_id_ld[29]) );
  AOI22_X1 U304 ( .A1(warp_checker_fence_regs_fence_en_ld[1]), .A2(n186), .B1(
        warp_gen_fence_regs_fence_en_ld[1]), .B2(n161), .ZN(n402) );
  AOI22_X1 U305 ( .A1(warp_checker_fence_regs_fence_en_ld[2]), .A2(n184), .B1(
        warp_gen_fence_regs_fence_en_ld[2]), .B2(n162), .ZN(n391) );
  AOI22_X1 U306 ( .A1(warp_checker_fence_regs_fence_en_ld[3]), .A2(n184), .B1(
        warp_gen_fence_regs_fence_en_ld[3]), .B2(n161), .ZN(n388) );
  AOI22_X1 U307 ( .A1(warp_checker_fence_regs_fence_en_ld[5]), .A2(n189), .B1(
        warp_gen_fence_regs_fence_en_ld[5]), .B2(n161), .ZN(n386) );
  AOI22_X1 U308 ( .A1(warp_checker_fence_regs_fence_en_ld[6]), .A2(n184), .B1(
        warp_gen_fence_regs_fence_en_ld[6]), .B2(n161), .ZN(n385) );
  AOI22_X1 U309 ( .A1(warp_checker_fence_regs_fence_en_ld[8]), .A2(n189), .B1(
        warp_gen_fence_regs_fence_en_ld[8]), .B2(n161), .ZN(n383) );
  AOI22_X1 U310 ( .A1(warp_checker_fence_regs_fence_en_ld[16]), .A2(n183), 
        .B1(warp_gen_fence_regs_fence_en_ld[16]), .B2(n162), .ZN(n406) );
  AOI22_X1 U311 ( .A1(warp_checker_fence_regs_fence_en_ld[17]), .A2(n186), 
        .B1(warp_gen_fence_regs_fence_en_ld[17]), .B2(n161), .ZN(n405) );
  AOI22_X1 U312 ( .A1(warp_checker_fence_regs_fence_en_ld[18]), .A2(n186), 
        .B1(warp_gen_fence_regs_fence_en_ld[18]), .B2(n162), .ZN(n404) );
  AOI22_X1 U313 ( .A1(warp_checker_fence_regs_fence_en_ld[19]), .A2(n183), 
        .B1(warp_gen_fence_regs_fence_en_ld[19]), .B2(n162), .ZN(n403) );
  AOI22_X1 U314 ( .A1(warp_checker_fence_regs_fence_en_ld[21]), .A2(n183), 
        .B1(warp_gen_fence_regs_fence_en_ld[21]), .B2(n162), .ZN(n400) );
  AOI22_X1 U315 ( .A1(warp_checker_fence_regs_fence_en_ld[22]), .A2(n187), 
        .B1(warp_gen_fence_regs_fence_en_ld[22]), .B2(n161), .ZN(n399) );
  AOI22_X1 U316 ( .A1(warp_checker_fence_regs_fence_en_ld[23]), .A2(n187), 
        .B1(warp_gen_fence_regs_fence_en_ld[23]), .B2(n162), .ZN(n398) );
  AOI22_X1 U317 ( .A1(warp_checker_fence_regs_fence_en_ld[24]), .A2(n183), 
        .B1(warp_gen_fence_regs_fence_en_ld[24]), .B2(n162), .ZN(n397) );
  AOI22_X1 U318 ( .A1(warp_checker_fence_regs_fence_en_ld[25]), .A2(n187), 
        .B1(warp_gen_fence_regs_fence_en_ld[25]), .B2(n161), .ZN(n396) );
  AOI22_X1 U319 ( .A1(warp_checker_fence_regs_fence_en_ld[26]), .A2(n188), 
        .B1(warp_gen_fence_regs_fence_en_ld[26]), .B2(n162), .ZN(n395) );
  AOI22_X1 U320 ( .A1(warp_checker_fence_regs_fence_en_ld[29]), .A2(n184), 
        .B1(warp_gen_fence_regs_fence_en_ld[29]), .B2(n162), .ZN(n392) );
  AOI22_X1 U321 ( .A1(warp_checker_fence_regs_fence_en_ld[31]), .A2(n188), 
        .B1(warp_gen_fence_regs_fence_en_ld[31]), .B2(n161), .ZN(n389) );
  AOI22_X1 U322 ( .A1(warp_checker_fence_regs_fence_en_ld[4]), .A2(n189), .B1(
        warp_gen_fence_regs_fence_en_ld[4]), .B2(n160), .ZN(n387) );
  AOI22_X1 U323 ( .A1(warp_checker_fence_regs_fence_en_ld[7]), .A2(n182), .B1(
        warp_gen_fence_regs_fence_en_ld[7]), .B2(n160), .ZN(n384) );
  AOI22_X1 U324 ( .A1(warp_checker_fence_regs_fence_en_ld[9]), .A2(n185), .B1(
        warp_gen_fence_regs_fence_en_ld[9]), .B2(n160), .ZN(n382) );
  AOI22_X1 U325 ( .A1(warp_checker_fence_regs_fence_en_ld[11]), .A2(n185), 
        .B1(warp_gen_fence_regs_fence_en_ld[11]), .B2(n160), .ZN(n411) );
  AOI22_X1 U326 ( .A1(warp_checker_fence_regs_fence_en_ld[14]), .A2(n182), 
        .B1(warp_gen_fence_regs_fence_en_ld[14]), .B2(n160), .ZN(n408) );
  AOI22_X1 U327 ( .A1(warp_checker_fence_regs_fence_en_ld[20]), .A2(n187), 
        .B1(warp_gen_fence_regs_fence_en_ld[20]), .B2(n160), .ZN(n401) );
  AOI22_X1 U328 ( .A1(warp_checker_fence_regs_fence_en_ld[27]), .A2(n182), 
        .B1(warp_gen_fence_regs_fence_en_ld[27]), .B2(n160), .ZN(n394) );
  AOI22_X1 U329 ( .A1(warp_checker_fence_regs_fence_en_ld[28]), .A2(n188), 
        .B1(warp_gen_fence_regs_fence_en_ld[28]), .B2(n160), .ZN(n393) );
  AOI22_X1 U330 ( .A1(warp_checker_fence_regs_fence_en_ld[30]), .A2(n188), 
        .B1(warp_gen_fence_regs_fence_en_ld[30]), .B2(n160), .ZN(n390) );
  AOI22_X1 U331 ( .A1(warp_checker_fence_regs_fence_en_ld[10]), .A2(n181), 
        .B1(warp_gen_fence_regs_fence_en_ld[10]), .B2(n163), .ZN(n412) );
  AOI22_X1 U332 ( .A1(warp_checker_fence_regs_fence_en_ld[12]), .A2(n185), 
        .B1(warp_gen_fence_regs_fence_en_ld[12]), .B2(n163), .ZN(n410) );
  AOI22_X1 U333 ( .A1(warp_checker_fence_regs_fence_en_ld[13]), .A2(n182), 
        .B1(warp_gen_fence_regs_fence_en_ld[13]), .B2(n163), .ZN(n409) );
  AOI22_X1 U334 ( .A1(warp_checker_fence_regs_fence_en_ld[15]), .A2(n186), 
        .B1(warp_gen_fence_regs_fence_en_ld[15]), .B2(n163), .ZN(n407) );
  AOI22_X1 U335 ( .A1(warp_checker_fence_regs_fence_en_ld[0]), .A2(n185), .B1(
        warp_gen_fence_regs_fence_en_ld[0]), .B2(n163), .ZN(n413) );
  AND2_X1 U336 ( .A1(\warp_gen_fence_regs_wr_cta_id[10><0] ), .A2(n173), .ZN(
        \fence_regs_wr_cta_id[10><0] ) );
  AND2_X1 U337 ( .A1(\warp_gen_fence_regs_wr_cta_id[11><0] ), .A2(n164), .ZN(
        \fence_regs_wr_cta_id[11><0] ) );
  AND2_X1 U338 ( .A1(\warp_gen_fence_regs_wr_cta_id[12><0] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[12><0] ) );
  AND2_X1 U339 ( .A1(\warp_gen_fence_regs_wr_cta_id[13><0] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[13><0] ) );
  AND2_X1 U340 ( .A1(\warp_gen_fence_regs_wr_cta_id[14><0] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[14><0] ) );
  AND2_X1 U341 ( .A1(\warp_gen_fence_regs_wr_cta_id[15><0] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[15><0] ) );
  AND2_X1 U342 ( .A1(\warp_gen_fence_regs_wr_cta_id[16><0] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[16><0] ) );
  AND2_X1 U343 ( .A1(\warp_gen_fence_regs_wr_cta_id[0><0] ), .A2(n173), .ZN(
        \fence_regs_wr_cta_id[0><0] ) );
  AND2_X1 U344 ( .A1(\warp_gen_fence_regs_wr_cta_id[1><0] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[1><0] ) );
  AND2_X1 U345 ( .A1(\warp_gen_fence_regs_wr_cta_id[2><0] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[2><0] ) );
  AND2_X1 U346 ( .A1(\warp_gen_fence_regs_wr_cta_id[17><0] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[17><0] ) );
  AND2_X1 U347 ( .A1(\warp_gen_fence_regs_wr_cta_id[18><0] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[18><0] ) );
  AND2_X1 U348 ( .A1(\warp_gen_fence_regs_wr_cta_id[19><0] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[19><0] ) );
  AND2_X1 U349 ( .A1(\warp_gen_fence_regs_wr_cta_id[20><0] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[20><0] ) );
  AND2_X1 U350 ( .A1(\warp_gen_fence_regs_wr_cta_id[21><0] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[21><0] ) );
  AND2_X1 U351 ( .A1(\warp_gen_fence_regs_wr_cta_id[22><0] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[22><0] ) );
  AND2_X1 U352 ( .A1(\warp_gen_fence_regs_wr_cta_id[23><0] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[23><0] ) );
  AND2_X1 U353 ( .A1(\warp_gen_fence_regs_wr_cta_id[24><0] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[24><0] ) );
  AND2_X1 U354 ( .A1(\warp_gen_fence_regs_wr_cta_id[25><0] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[25><0] ) );
  AND2_X1 U355 ( .A1(\warp_gen_fence_regs_wr_cta_id[26><0] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[26><0] ) );
  AND2_X1 U356 ( .A1(\warp_gen_fence_regs_wr_cta_id[27><0] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[27><0] ) );
  AND2_X1 U357 ( .A1(\warp_gen_fence_regs_wr_cta_id[28><0] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[28><0] ) );
  AND2_X1 U358 ( .A1(\warp_gen_fence_regs_wr_cta_id[29><0] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[29><0] ) );
  AND2_X1 U359 ( .A1(\warp_gen_fence_regs_wr_cta_id[10><1] ), .A2(n173), .ZN(
        \fence_regs_wr_cta_id[10><1] ) );
  AND2_X1 U360 ( .A1(\warp_gen_fence_regs_wr_cta_id[10><2] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[10><2] ) );
  AND2_X1 U361 ( .A1(\warp_gen_fence_regs_wr_cta_id[10><3] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[10><3] ) );
  AND2_X1 U362 ( .A1(\warp_gen_fence_regs_wr_cta_id[11><1] ), .A2(n164), .ZN(
        \fence_regs_wr_cta_id[11><1] ) );
  AND2_X1 U363 ( .A1(\warp_gen_fence_regs_wr_cta_id[11><2] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[11><2] ) );
  AND2_X1 U364 ( .A1(\warp_gen_fence_regs_wr_cta_id[11><3] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[11><3] ) );
  AND2_X1 U365 ( .A1(\warp_gen_fence_regs_wr_cta_id[12><1] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[12><1] ) );
  AND2_X1 U366 ( .A1(\warp_gen_fence_regs_wr_cta_id[12><2] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[12><2] ) );
  AND2_X1 U367 ( .A1(\warp_gen_fence_regs_wr_cta_id[12><3] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[12><3] ) );
  AND2_X1 U368 ( .A1(\warp_gen_fence_regs_wr_cta_id[13><1] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[13><1] ) );
  AND2_X1 U369 ( .A1(\warp_gen_fence_regs_wr_cta_id[13><2] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[13><2] ) );
  AND2_X1 U370 ( .A1(\warp_gen_fence_regs_wr_cta_id[13><3] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[13><3] ) );
  AND2_X1 U371 ( .A1(\warp_gen_fence_regs_wr_cta_id[14><1] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[14><1] ) );
  AND2_X1 U372 ( .A1(\warp_gen_fence_regs_wr_cta_id[14><2] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[14><2] ) );
  AND2_X1 U373 ( .A1(\warp_gen_fence_regs_wr_cta_id[14><3] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[14><3] ) );
  AND2_X1 U374 ( .A1(\warp_gen_fence_regs_wr_cta_id[15><1] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[15><1] ) );
  AND2_X1 U375 ( .A1(\warp_gen_fence_regs_wr_cta_id[15><2] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[15><2] ) );
  AND2_X1 U376 ( .A1(\warp_gen_fence_regs_wr_cta_id[15><3] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[15><3] ) );
  AND2_X1 U377 ( .A1(\warp_gen_fence_regs_wr_cta_id[16><1] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[16><1] ) );
  AND2_X1 U378 ( .A1(\warp_gen_fence_regs_wr_cta_id[16><2] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[16><2] ) );
  AND2_X1 U379 ( .A1(\warp_gen_fence_regs_wr_cta_id[16><3] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[16><3] ) );
  AND2_X1 U380 ( .A1(\warp_gen_fence_regs_wr_cta_id[0><1] ), .A2(n173), .ZN(
        \fence_regs_wr_cta_id[0><1] ) );
  AND2_X1 U381 ( .A1(\warp_gen_fence_regs_wr_cta_id[0><2] ), .A2(n173), .ZN(
        \fence_regs_wr_cta_id[0><2] ) );
  AND2_X1 U382 ( .A1(\warp_gen_fence_regs_wr_cta_id[0><3] ), .A2(n173), .ZN(
        \fence_regs_wr_cta_id[0><3] ) );
  AND2_X1 U383 ( .A1(\warp_gen_fence_regs_wr_cta_id[1><1] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[1><1] ) );
  AND2_X1 U384 ( .A1(\warp_gen_fence_regs_wr_cta_id[1><2] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[1><2] ) );
  AND2_X1 U385 ( .A1(\warp_gen_fence_regs_wr_cta_id[1><3] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[1><3] ) );
  AND2_X1 U386 ( .A1(\warp_gen_fence_regs_wr_cta_id[2><1] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[2><1] ) );
  AND2_X1 U387 ( .A1(\warp_gen_fence_regs_wr_cta_id[2><2] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[2><2] ) );
  AND2_X1 U388 ( .A1(\warp_gen_fence_regs_wr_cta_id[2><3] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[2><3] ) );
  AND2_X1 U389 ( .A1(\warp_gen_fence_regs_wr_cta_id[17><1] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[17><1] ) );
  AND2_X1 U390 ( .A1(\warp_gen_fence_regs_wr_cta_id[17><2] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[17><2] ) );
  AND2_X1 U391 ( .A1(\warp_gen_fence_regs_wr_cta_id[17><3] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[17><3] ) );
  AND2_X1 U392 ( .A1(\warp_gen_fence_regs_wr_cta_id[18><1] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[18><1] ) );
  AND2_X1 U393 ( .A1(\warp_gen_fence_regs_wr_cta_id[18><2] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[18><2] ) );
  AND2_X1 U394 ( .A1(\warp_gen_fence_regs_wr_cta_id[18><3] ), .A2(n166), .ZN(
        \fence_regs_wr_cta_id[18><3] ) );
  AND2_X1 U395 ( .A1(\warp_gen_fence_regs_wr_cta_id[19><1] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[19><1] ) );
  AND2_X1 U396 ( .A1(\warp_gen_fence_regs_wr_cta_id[19><2] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[19><2] ) );
  AND2_X1 U397 ( .A1(\warp_gen_fence_regs_wr_cta_id[19><3] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[19><3] ) );
  AND2_X1 U398 ( .A1(\warp_gen_fence_regs_wr_cta_id[20><1] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[20><1] ) );
  AND2_X1 U399 ( .A1(\warp_gen_fence_regs_wr_cta_id[20><2] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[20><2] ) );
  AND2_X1 U400 ( .A1(\warp_gen_fence_regs_wr_cta_id[20><3] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[20><3] ) );
  AND2_X1 U401 ( .A1(\warp_gen_fence_regs_wr_cta_id[21><1] ), .A2(n167), .ZN(
        \fence_regs_wr_cta_id[21><1] ) );
  AND2_X1 U402 ( .A1(\warp_gen_fence_regs_wr_cta_id[21><2] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[21><2] ) );
  AND2_X1 U403 ( .A1(\warp_gen_fence_regs_wr_cta_id[21><3] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[21><3] ) );
  AND2_X1 U404 ( .A1(\warp_gen_fence_regs_wr_cta_id[22><1] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[22><1] ) );
  AND2_X1 U405 ( .A1(\warp_gen_fence_regs_wr_cta_id[22><2] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[22><2] ) );
  AND2_X1 U406 ( .A1(\warp_gen_fence_regs_wr_cta_id[22><3] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[22><3] ) );
  AND2_X1 U407 ( .A1(\warp_gen_fence_regs_wr_cta_id[23><1] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[23><1] ) );
  AND2_X1 U408 ( .A1(\warp_gen_fence_regs_wr_cta_id[23><2] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[23><2] ) );
  AND2_X1 U409 ( .A1(\warp_gen_fence_regs_wr_cta_id[23><3] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[23><3] ) );
  AND2_X1 U410 ( .A1(\warp_gen_fence_regs_wr_cta_id[24><1] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[24><1] ) );
  AND2_X1 U411 ( .A1(\warp_gen_fence_regs_wr_cta_id[24><2] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[24><2] ) );
  AND2_X1 U412 ( .A1(\warp_gen_fence_regs_wr_cta_id[24><3] ), .A2(n168), .ZN(
        \fence_regs_wr_cta_id[24><3] ) );
  AND2_X1 U413 ( .A1(\warp_gen_fence_regs_wr_cta_id[25><1] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[25><1] ) );
  AND2_X1 U414 ( .A1(\warp_gen_fence_regs_wr_cta_id[25><2] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[25><2] ) );
  AND2_X1 U415 ( .A1(\warp_gen_fence_regs_wr_cta_id[25><3] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[25><3] ) );
  AND2_X1 U416 ( .A1(\warp_gen_fence_regs_wr_cta_id[26><1] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[26><1] ) );
  AND2_X1 U417 ( .A1(\warp_gen_fence_regs_wr_cta_id[26><2] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[26><2] ) );
  AND2_X1 U418 ( .A1(\warp_gen_fence_regs_wr_cta_id[26><3] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[26><3] ) );
  AND2_X1 U419 ( .A1(\warp_gen_fence_regs_wr_cta_id[27><1] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[27><1] ) );
  AND2_X1 U420 ( .A1(\warp_gen_fence_regs_wr_cta_id[27><2] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[27><2] ) );
  AND2_X1 U421 ( .A1(\warp_gen_fence_regs_wr_cta_id[27><3] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[27><3] ) );
  AND2_X1 U422 ( .A1(\warp_gen_fence_regs_wr_cta_id[28><1] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[28><1] ) );
  AND2_X1 U423 ( .A1(\warp_gen_fence_regs_wr_cta_id[28><2] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[28><2] ) );
  AND2_X1 U424 ( .A1(\warp_gen_fence_regs_wr_cta_id[28><3] ), .A2(n169), .ZN(
        \fence_regs_wr_cta_id[28><3] ) );
  AND2_X1 U425 ( .A1(\warp_gen_fence_regs_wr_cta_id[29><1] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[29><1] ) );
  AND2_X1 U426 ( .A1(\warp_gen_fence_regs_wr_cta_id[29><2] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[29><2] ) );
  AND2_X1 U427 ( .A1(\warp_gen_fence_regs_wr_cta_id[29><3] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[29><3] ) );
  INV_X1 U428 ( .A(n387), .ZN(n5) );
  INV_X1 U429 ( .A(n384), .ZN(n8) );
  INV_X1 U430 ( .A(n382), .ZN(n10) );
  INV_X1 U431 ( .A(n411), .ZN(n12) );
  INV_X1 U432 ( .A(n408), .ZN(n15) );
  INV_X1 U433 ( .A(n401), .ZN(n21) );
  INV_X1 U434 ( .A(n394), .ZN(n28) );
  INV_X1 U435 ( .A(n393), .ZN(n29) );
  INV_X1 U436 ( .A(n390), .ZN(n31) );
  AND2_X1 U437 ( .A1(\warp_gen_fence_regs_wr_cta_id[3><0] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[3><0] ) );
  AND2_X1 U438 ( .A1(\warp_gen_fence_regs_wr_cta_id[3><1] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[3><1] ) );
  AND2_X1 U439 ( .A1(\warp_gen_fence_regs_wr_cta_id[3><2] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[3><2] ) );
  AND2_X1 U440 ( .A1(\warp_gen_fence_regs_wr_cta_id[3><3] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[3><3] ) );
  AND2_X1 U441 ( .A1(\warp_gen_fence_regs_wr_cta_id[4><0] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[4><0] ) );
  AND2_X1 U442 ( .A1(\warp_gen_fence_regs_wr_cta_id[4><1] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[4><1] ) );
  AND2_X1 U443 ( .A1(\warp_gen_fence_regs_wr_cta_id[4><2] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[4><2] ) );
  AND2_X1 U444 ( .A1(\warp_gen_fence_regs_wr_cta_id[4><3] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[4><3] ) );
  AND2_X1 U445 ( .A1(\warp_gen_fence_regs_wr_cta_id[5><0] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[5><0] ) );
  AND2_X1 U446 ( .A1(\warp_gen_fence_regs_wr_cta_id[5><1] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[5><1] ) );
  AND2_X1 U447 ( .A1(\warp_gen_fence_regs_wr_cta_id[5><2] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[5><2] ) );
  AND2_X1 U448 ( .A1(\warp_gen_fence_regs_wr_cta_id[5><3] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[5><3] ) );
  AND2_X1 U449 ( .A1(\warp_gen_fence_regs_wr_cta_id[6><0] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[6><0] ) );
  AND2_X1 U450 ( .A1(\warp_gen_fence_regs_wr_cta_id[6><1] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[6><1] ) );
  AND2_X1 U451 ( .A1(\warp_gen_fence_regs_wr_cta_id[6><2] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[6><2] ) );
  AND2_X1 U452 ( .A1(\warp_gen_fence_regs_wr_cta_id[6><3] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[6><3] ) );
  AND2_X1 U453 ( .A1(\warp_gen_fence_regs_wr_cta_id[7><0] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[7><0] ) );
  AND2_X1 U454 ( .A1(\warp_gen_fence_regs_wr_cta_id[7><1] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[7><1] ) );
  AND2_X1 U455 ( .A1(\warp_gen_fence_regs_wr_cta_id[7><2] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[7><2] ) );
  AND2_X1 U456 ( .A1(\warp_gen_fence_regs_wr_cta_id[7><3] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[7><3] ) );
  AND2_X1 U457 ( .A1(\warp_gen_fence_regs_wr_cta_id[8><0] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[8><0] ) );
  AND2_X1 U458 ( .A1(\warp_gen_fence_regs_wr_cta_id[8><1] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[8><1] ) );
  AND2_X1 U459 ( .A1(\warp_gen_fence_regs_wr_cta_id[8><2] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[8><2] ) );
  AND2_X1 U460 ( .A1(\warp_gen_fence_regs_wr_cta_id[8><3] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[8><3] ) );
  AND2_X1 U461 ( .A1(\warp_gen_fence_regs_wr_cta_id[9><0] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[9><0] ) );
  AND2_X1 U462 ( .A1(\warp_gen_fence_regs_wr_cta_id[9><1] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[9><1] ) );
  AND2_X1 U463 ( .A1(\warp_gen_fence_regs_wr_cta_id[9><2] ), .A2(n172), .ZN(
        \fence_regs_wr_cta_id[9><2] ) );
  AND2_X1 U464 ( .A1(\warp_gen_fence_regs_wr_cta_id[9><3] ), .A2(n165), .ZN(
        \fence_regs_wr_cta_id[9><3] ) );
  AND2_X1 U465 ( .A1(\warp_gen_fence_regs_wr_cta_id[30><0] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[30><0] ) );
  AND2_X1 U466 ( .A1(\warp_gen_fence_regs_wr_cta_id[30><1] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[30><1] ) );
  AND2_X1 U467 ( .A1(\warp_gen_fence_regs_wr_cta_id[30><2] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[30><2] ) );
  AND2_X1 U468 ( .A1(\warp_gen_fence_regs_wr_cta_id[30><3] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[30><3] ) );
  AND2_X1 U469 ( .A1(\warp_gen_fence_regs_wr_cta_id[31><0] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[31><0] ) );
  AND2_X1 U470 ( .A1(\warp_gen_fence_regs_wr_cta_id[31><1] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[31><1] ) );
  AND2_X1 U471 ( .A1(\warp_gen_fence_regs_wr_cta_id[31><2] ), .A2(n170), .ZN(
        \fence_regs_wr_cta_id[31><2] ) );
  AND2_X1 U472 ( .A1(\warp_gen_fence_regs_wr_cta_id[31><3] ), .A2(n171), .ZN(
        \fence_regs_wr_cta_id[31><3] ) );
  INV_X1 U473 ( .A(n402), .ZN(n2) );
  INV_X1 U474 ( .A(n391), .ZN(n3) );
  INV_X1 U475 ( .A(n388), .ZN(n4) );
  INV_X1 U476 ( .A(n386), .ZN(n6) );
  INV_X1 U477 ( .A(n385), .ZN(n7) );
  INV_X1 U478 ( .A(n383), .ZN(n9) );
  INV_X1 U479 ( .A(n406), .ZN(n17) );
  INV_X1 U480 ( .A(n405), .ZN(n18) );
  INV_X1 U481 ( .A(n404), .ZN(n19) );
  INV_X1 U482 ( .A(n403), .ZN(n20) );
  INV_X1 U483 ( .A(n400), .ZN(n22) );
  INV_X1 U484 ( .A(n399), .ZN(n23) );
  INV_X1 U485 ( .A(n398), .ZN(n24) );
  INV_X1 U486 ( .A(n397), .ZN(n25) );
  INV_X1 U487 ( .A(n396), .ZN(n26) );
  INV_X1 U488 ( .A(n395), .ZN(n27) );
  INV_X1 U489 ( .A(n392), .ZN(n30) );
  INV_X1 U490 ( .A(n389), .ZN(n32) );
  INV_X1 U491 ( .A(n412), .ZN(n11) );
  INV_X1 U492 ( .A(n410), .ZN(n13) );
  INV_X1 U493 ( .A(n409), .ZN(n14) );
  INV_X1 U494 ( .A(n407), .ZN(n16) );
  INV_X1 U495 ( .A(n413), .ZN(n1) );
  BUF_X1 U496 ( .A(host_reset), .Z(n248) );
  BUF_X1 U497 ( .A(host_reset), .Z(n249) );
  AND2_X1 U498 ( .A1(warp_gen_pool_wr_data[101]), .A2(n176), .ZN(n65) );
  AND2_X1 U499 ( .A1(warp_gen_pool_wr_data[102]), .A2(n176), .ZN(n66) );
  AND2_X1 U500 ( .A1(warp_gen_pool_wr_data[103]), .A2(n176), .ZN(n67) );
  AND2_X1 U501 ( .A1(warp_gen_pool_wr_data[104]), .A2(n176), .ZN(n68) );
  AND2_X1 U502 ( .A1(warp_gen_pool_wr_data[105]), .A2(n176), .ZN(n69) );
  AND2_X1 U503 ( .A1(warp_gen_pool_wr_data[106]), .A2(n176), .ZN(n70) );
  AND2_X1 U504 ( .A1(warp_gen_pool_wr_data[107]), .A2(n176), .ZN(n71) );
  AND2_X1 U505 ( .A1(warp_gen_pool_wr_data[108]), .A2(n176), .ZN(n72) );
  AND2_X1 U506 ( .A1(warp_gen_pool_wr_data[109]), .A2(n176), .ZN(n73) );
  AND2_X1 U507 ( .A1(warp_gen_pool_wr_data[110]), .A2(n176), .ZN(n74) );
  AND2_X1 U508 ( .A1(warp_gen_pool_wr_data[111]), .A2(n176), .ZN(n75) );
  AND2_X1 U509 ( .A1(warp_gen_pool_wr_data[112]), .A2(n176), .ZN(n76) );
  AND2_X1 U510 ( .A1(warp_gen_pool_wr_data[113]), .A2(n176), .ZN(n77) );
  AND2_X1 U511 ( .A1(warp_gen_pool_wr_data[114]), .A2(n176), .ZN(n78) );
  AND2_X1 U512 ( .A1(warp_gen_pool_wr_data[115]), .A2(n176), .ZN(n79) );
  AND2_X1 U513 ( .A1(warp_gen_pool_wr_data[116]), .A2(n176), .ZN(n80) );
  INV_X1 U514 ( .A(n208), .ZN(n251) );
  AOI22_X1 U515 ( .A1(n164), .A2(warp_gen_state_wr_en), .B1(
        warp_sched_state_wr_en), .B2(n181), .ZN(n208) );
  INV_X1 U516 ( .A(n214), .ZN(n260) );
  AOI22_X1 U517 ( .A1(warp_gen_state_addr[1]), .A2(n163), .B1(
        warp_sched_state_addr[1]), .B2(n179), .ZN(n214) );
  INV_X1 U518 ( .A(n213), .ZN(n254) );
  AOI22_X1 U519 ( .A1(warp_gen_state_addr[2]), .A2(n163), .B1(
        warp_sched_state_addr[2]), .B2(n179), .ZN(n213) );
  INV_X1 U520 ( .A(n346), .ZN(n253) );
  AOI22_X1 U521 ( .A1(warp_gen_pool_addr[3]), .A2(n163), .B1(
        warp_sched_pool_addr[3]), .B2(n180), .ZN(n346) );
  INV_X1 U522 ( .A(n345), .ZN(n259) );
  AOI22_X1 U523 ( .A1(warp_gen_pool_addr[4]), .A2(n163), .B1(
        warp_sched_pool_addr[4]), .B2(n180), .ZN(n345) );
  INV_X1 U524 ( .A(n215), .ZN(n256) );
  AOI22_X1 U525 ( .A1(warp_gen_state_addr[0]), .A2(n164), .B1(
        warp_sched_state_addr[0]), .B2(n180), .ZN(n215) );
  INV_X1 U526 ( .A(n212), .ZN(n252) );
  AOI22_X1 U527 ( .A1(warp_gen_state_addr[3]), .A2(n164), .B1(
        warp_sched_state_addr[3]), .B2(n179), .ZN(n212) );
  INV_X1 U528 ( .A(n211), .ZN(n258) );
  AOI22_X1 U529 ( .A1(warp_gen_state_addr[4]), .A2(n164), .B1(
        warp_sched_state_addr[4]), .B2(n179), .ZN(n211) );
  INV_X1 U530 ( .A(n349), .ZN(n257) );
  AOI22_X1 U531 ( .A1(warp_gen_pool_addr[0]), .A2(n164), .B1(
        warp_sched_pool_addr[0]), .B2(n181), .ZN(n349) );
  INV_X1 U532 ( .A(n348), .ZN(n261) );
  AOI22_X1 U533 ( .A1(warp_gen_pool_addr[1]), .A2(n164), .B1(
        warp_sched_pool_addr[1]), .B2(n181), .ZN(n348) );
  INV_X1 U534 ( .A(n347), .ZN(n255) );
  AOI22_X1 U535 ( .A1(warp_gen_pool_addr[2]), .A2(n164), .B1(
        warp_sched_pool_addr[2]), .B2(n180), .ZN(n347) );
  AND2_X1 U536 ( .A1(warp_gen_pool_wr_data[0]), .A2(n175), .ZN(n81) );
  AND2_X1 U537 ( .A1(warp_gen_pool_wr_data[117]), .A2(n175), .ZN(n82) );
  AND2_X1 U538 ( .A1(warp_gen_pool_wr_data[118]), .A2(n175), .ZN(n83) );
  AND2_X1 U539 ( .A1(warp_gen_pool_wr_data[119]), .A2(n175), .ZN(n84) );
  AND2_X1 U540 ( .A1(warp_gen_pool_wr_data[120]), .A2(n175), .ZN(n85) );
  AND2_X1 U541 ( .A1(warp_gen_pool_wr_data[121]), .A2(n175), .ZN(n86) );
  AND2_X1 U542 ( .A1(warp_gen_pool_wr_data[122]), .A2(n175), .ZN(n87) );
  AND2_X1 U543 ( .A1(warp_gen_pool_wr_data[123]), .A2(n175), .ZN(n88) );
  AND2_X1 U544 ( .A1(warp_gen_pool_wr_en), .A2(n178), .ZN(n89) );
  AND2_X1 U545 ( .A1(warp_gen_pool_wr_data[37]), .A2(n177), .ZN(n90) );
  AND2_X1 U546 ( .A1(warp_gen_pool_wr_data[38]), .A2(n178), .ZN(n91) );
  AND2_X1 U547 ( .A1(warp_gen_pool_wr_data[39]), .A2(n176), .ZN(n92) );
  AND2_X1 U548 ( .A1(warp_gen_pool_wr_data[40]), .A2(n178), .ZN(n93) );
  AND2_X1 U549 ( .A1(warp_gen_pool_wr_data[41]), .A2(n177), .ZN(n94) );
  AND2_X1 U550 ( .A1(warp_gen_pool_wr_data[42]), .A2(n177), .ZN(n95) );
  AND2_X1 U551 ( .A1(warp_gen_pool_wr_data[43]), .A2(n176), .ZN(n96) );
  AND2_X1 U552 ( .A1(warp_gen_pool_wr_data[44]), .A2(n178), .ZN(n97) );
  AND2_X1 U553 ( .A1(warp_gen_pool_wr_data[45]), .A2(n177), .ZN(n98) );
  AND2_X1 U554 ( .A1(warp_gen_pool_wr_data[46]), .A2(n176), .ZN(n99) );
  AND2_X1 U555 ( .A1(warp_gen_pool_wr_data[47]), .A2(n176), .ZN(n100) );
  AND2_X1 U556 ( .A1(warp_gen_pool_wr_data[48]), .A2(n178), .ZN(n101) );
  AND2_X1 U557 ( .A1(warp_gen_pool_wr_data[49]), .A2(n177), .ZN(n102) );
  AND2_X1 U558 ( .A1(warp_gen_pool_wr_data[50]), .A2(n178), .ZN(n103) );
  AND2_X1 U559 ( .A1(warp_gen_pool_wr_data[51]), .A2(n176), .ZN(n104) );
  AND2_X1 U560 ( .A1(warp_gen_pool_wr_data[5]), .A2(n178), .ZN(n105) );
  AND2_X1 U561 ( .A1(warp_gen_pool_wr_data[6]), .A2(n178), .ZN(n106) );
  AND2_X1 U562 ( .A1(warp_gen_pool_wr_data[7]), .A2(n178), .ZN(n107) );
  AND2_X1 U563 ( .A1(warp_gen_pool_wr_data[8]), .A2(n178), .ZN(n108) );
  AND2_X1 U564 ( .A1(warp_gen_pool_wr_data[9]), .A2(n178), .ZN(n109) );
  AND2_X1 U565 ( .A1(warp_gen_pool_wr_data[10]), .A2(n178), .ZN(n110) );
  AND2_X1 U566 ( .A1(warp_gen_pool_wr_data[11]), .A2(n178), .ZN(n111) );
  AND2_X1 U567 ( .A1(warp_gen_pool_wr_data[12]), .A2(n178), .ZN(n112) );
  AND2_X1 U568 ( .A1(warp_gen_pool_wr_data[13]), .A2(n178), .ZN(n113) );
  AND2_X1 U569 ( .A1(warp_gen_pool_wr_data[14]), .A2(n178), .ZN(n114) );
  AND2_X1 U570 ( .A1(warp_gen_pool_wr_data[15]), .A2(n178), .ZN(n115) );
  AND2_X1 U571 ( .A1(warp_gen_pool_wr_data[16]), .A2(n178), .ZN(n116) );
  AND2_X1 U572 ( .A1(warp_gen_pool_wr_data[17]), .A2(n178), .ZN(n117) );
  AND2_X1 U573 ( .A1(warp_gen_pool_wr_data[18]), .A2(n178), .ZN(n118) );
  AND2_X1 U574 ( .A1(warp_gen_pool_wr_data[19]), .A2(n178), .ZN(n119) );
  AND2_X1 U575 ( .A1(warp_gen_pool_wr_data[20]), .A2(n178), .ZN(n120) );
  AND2_X1 U576 ( .A1(warp_gen_pool_wr_data[21]), .A2(n177), .ZN(n121) );
  AND2_X1 U577 ( .A1(warp_gen_pool_wr_data[22]), .A2(n177), .ZN(n122) );
  AND2_X1 U578 ( .A1(warp_gen_pool_wr_data[23]), .A2(n177), .ZN(n123) );
  AND2_X1 U579 ( .A1(warp_gen_pool_wr_data[24]), .A2(n177), .ZN(n124) );
  AND2_X1 U580 ( .A1(warp_gen_pool_wr_data[25]), .A2(n177), .ZN(n125) );
  AND2_X1 U581 ( .A1(warp_gen_pool_wr_data[26]), .A2(n177), .ZN(n126) );
  AND2_X1 U582 ( .A1(warp_gen_pool_wr_data[27]), .A2(n177), .ZN(n127) );
  AND2_X1 U583 ( .A1(warp_gen_pool_wr_data[28]), .A2(n177), .ZN(n128) );
  AND2_X1 U584 ( .A1(warp_gen_pool_wr_data[29]), .A2(n177), .ZN(n129) );
  AND2_X1 U585 ( .A1(warp_gen_pool_wr_data[30]), .A2(n177), .ZN(n130) );
  AND2_X1 U586 ( .A1(warp_gen_pool_wr_data[31]), .A2(n177), .ZN(n131) );
  AND2_X1 U587 ( .A1(warp_gen_pool_wr_data[32]), .A2(n177), .ZN(n132) );
  AND2_X1 U588 ( .A1(warp_gen_pool_wr_data[33]), .A2(n177), .ZN(n133) );
  AND2_X1 U589 ( .A1(warp_gen_pool_wr_data[34]), .A2(n177), .ZN(n134) );
  AND2_X1 U590 ( .A1(warp_gen_pool_wr_data[35]), .A2(n177), .ZN(n135) );
  AND2_X1 U591 ( .A1(warp_gen_pool_wr_data[36]), .A2(n177), .ZN(n136) );
  AND2_X1 U592 ( .A1(warp_gen_pool_wr_data[52]), .A2(n176), .ZN(n137) );
  AND2_X1 U593 ( .A1(warp_gen_pool_wr_data[53]), .A2(n178), .ZN(n138) );
  AND2_X1 U594 ( .A1(warp_gen_pool_wr_data[54]), .A2(n177), .ZN(n139) );
  AND2_X1 U595 ( .A1(warp_gen_pool_wr_data[55]), .A2(n176), .ZN(n140) );
  AND2_X1 U596 ( .A1(warp_gen_pool_wr_data[56]), .A2(n178), .ZN(n141) );
  AND2_X1 U597 ( .A1(warp_gen_pool_wr_data[57]), .A2(n177), .ZN(n142) );
  AND2_X1 U598 ( .A1(warp_gen_pool_wr_data[58]), .A2(n176), .ZN(n143) );
  AND2_X1 U599 ( .A1(warp_gen_pool_wr_data[59]), .A2(n178), .ZN(n144) );
  AND2_X1 U600 ( .A1(warp_gen_pool_wr_data[60]), .A2(n177), .ZN(n145) );
  AND2_X1 U601 ( .A1(warp_gen_pool_wr_data[61]), .A2(n176), .ZN(n146) );
  AND2_X1 U602 ( .A1(warp_gen_pool_wr_data[62]), .A2(n178), .ZN(n147) );
  AND2_X1 U603 ( .A1(warp_gen_pool_wr_data[63]), .A2(n177), .ZN(n148) );
  AND2_X1 U604 ( .A1(warp_gen_pool_wr_data[97]), .A2(n176), .ZN(n149) );
  AND2_X1 U605 ( .A1(warp_gen_pool_wr_data[98]), .A2(n178), .ZN(n150) );
  AND2_X1 U606 ( .A1(warp_gen_pool_wr_data[99]), .A2(n177), .ZN(n151) );
  AND2_X1 U607 ( .A1(warp_gen_pool_wr_data[100]), .A2(n176), .ZN(n152) );
  AND2_X1 U608 ( .A1(warp_gen_pool_wr_data[1]), .A2(n178), .ZN(n153) );
  AND2_X1 U609 ( .A1(warp_gen_pool_wr_data[2]), .A2(n177), .ZN(n154) );
  AND2_X1 U610 ( .A1(warp_gen_pool_wr_data[3]), .A2(n177), .ZN(n155) );
  AND2_X1 U611 ( .A1(warp_gen_pool_wr_data[4]), .A2(n176), .ZN(n156) );
  AND2_X1 U612 ( .A1(\warp_sched_state_wr_data[0] ), .A2(n224), .ZN(n157) );
  INV_X1 U613 ( .A(n220), .ZN(n161) );
  INV_X1 U614 ( .A(n220), .ZN(n162) );
  INV_X1 U615 ( .A(n219), .ZN(n166) );
  INV_X1 U616 ( .A(n220), .ZN(n168) );
  INV_X1 U617 ( .A(n219), .ZN(n169) );
  INV_X1 U618 ( .A(n221), .ZN(n173) );
  INV_X1 U619 ( .A(n221), .ZN(n176) );
endmodule
