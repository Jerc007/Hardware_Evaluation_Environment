


module warp_generator_SHMEM_ADDR_SIZE14_DW01_inc_1 ( A, SUM );
  input [11:0] A;
  output [11:0] SUM;

  wire   [11:2] carry;

  HA_X1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  HA_X1 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  HA_X1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(carry[11]), .B(A[11]), .Z(SUM[11]) );
  INV_X1 U2 ( .A(A[0]), .ZN(SUM[0]) );
endmodule


module warp_generator_SHMEM_ADDR_SIZE14_DW01_add_1 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46;

  OR2_X1 U2 ( .A1(B[3]), .A2(A[3]), .ZN(n1) );
  INV_X1 U3 ( .A(n19), .ZN(n7) );
  INV_X1 U4 ( .A(n41), .ZN(n5) );
  INV_X1 U5 ( .A(n28), .ZN(n10) );
  INV_X1 U6 ( .A(n44), .ZN(n8) );
  INV_X1 U7 ( .A(n35), .ZN(n11) );
  INV_X1 U8 ( .A(n30), .ZN(n9) );
  INV_X1 U9 ( .A(A[2]), .ZN(n12) );
  INV_X1 U10 ( .A(n16), .ZN(n6) );
  AND2_X1 U11 ( .A1(n36), .A2(n1), .ZN(SUM[3]) );
  BUF_X1 U12 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  XOR2_X1 U14 ( .A(n13), .B(n14), .Z(SUM[9]) );
  NAND2_X1 U15 ( .A1(n15), .A2(n6), .ZN(n13) );
  XOR2_X1 U16 ( .A(n17), .B(n18), .Z(SUM[8]) );
  NOR2_X1 U17 ( .A1(n19), .A2(n20), .ZN(n18) );
  XNOR2_X1 U18 ( .A(n21), .B(n22), .ZN(SUM[7]) );
  AND2_X1 U19 ( .A1(n23), .A2(n8), .ZN(n22) );
  AOI21_X1 U20 ( .B1(n24), .B2(n25), .A(n9), .ZN(n21) );
  XNOR2_X1 U21 ( .A(n26), .B(n24), .ZN(SUM[6]) );
  OAI21_X1 U22 ( .B1(n27), .B2(n28), .A(n29), .ZN(n24) );
  NAND2_X1 U23 ( .A1(n25), .A2(n30), .ZN(n26) );
  XNOR2_X1 U24 ( .A(n27), .B(n31), .ZN(SUM[5]) );
  AND2_X1 U25 ( .A1(n29), .A2(n10), .ZN(n31) );
  NOR2_X1 U26 ( .A1(n32), .A2(n11), .ZN(n27) );
  XNOR2_X1 U27 ( .A(n36), .B(n33), .ZN(SUM[4]) );
  NOR2_X1 U28 ( .A1(n34), .A2(n11), .ZN(n33) );
  INV_X1 U29 ( .A(n12), .ZN(SUM[2]) );
  XOR2_X1 U30 ( .A(n37), .B(n38), .Z(SUM[11]) );
  AOI21_X1 U31 ( .B1(n39), .B2(n5), .A(n40), .ZN(n38) );
  XNOR2_X1 U32 ( .A(B[11]), .B(A[11]), .ZN(n37) );
  XOR2_X1 U33 ( .A(n39), .B(n42), .Z(SUM[10]) );
  NOR2_X1 U34 ( .A1(n41), .A2(n40), .ZN(n42) );
  AND2_X1 U35 ( .A1(B[10]), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U36 ( .A1(B[10]), .A2(A[10]), .ZN(n41) );
  OAI21_X1 U37 ( .B1(n16), .B2(n14), .A(n15), .ZN(n39) );
  NAND2_X1 U38 ( .A1(B[9]), .A2(A[9]), .ZN(n15) );
  AOI21_X1 U39 ( .B1(n7), .B2(n17), .A(n20), .ZN(n14) );
  AND2_X1 U40 ( .A1(B[8]), .A2(A[8]), .ZN(n20) );
  OAI211_X1 U41 ( .C1(n43), .C2(n44), .A(n23), .B(n45), .ZN(n17) );
  NAND4_X1 U42 ( .A1(n32), .A2(n10), .A3(n25), .A4(n8), .ZN(n45) );
  NOR2_X1 U43 ( .A1(n36), .A2(n34), .ZN(n32) );
  NOR2_X1 U44 ( .A1(B[4]), .A2(A[4]), .ZN(n34) );
  NAND2_X1 U45 ( .A1(B[3]), .A2(A[3]), .ZN(n36) );
  NAND2_X1 U46 ( .A1(B[7]), .A2(A[7]), .ZN(n23) );
  NOR2_X1 U47 ( .A1(B[7]), .A2(A[7]), .ZN(n44) );
  AOI21_X1 U48 ( .B1(n25), .B2(n46), .A(n9), .ZN(n43) );
  NAND2_X1 U49 ( .A1(B[6]), .A2(A[6]), .ZN(n30) );
  OAI21_X1 U50 ( .B1(n28), .B2(n35), .A(n29), .ZN(n46) );
  NAND2_X1 U51 ( .A1(B[5]), .A2(A[5]), .ZN(n29) );
  NAND2_X1 U52 ( .A1(B[4]), .A2(A[4]), .ZN(n35) );
  NOR2_X1 U53 ( .A1(B[5]), .A2(A[5]), .ZN(n28) );
  OR2_X1 U54 ( .A1(B[6]), .A2(A[6]), .ZN(n25) );
  NOR2_X1 U55 ( .A1(B[8]), .A2(A[8]), .ZN(n19) );
  NOR2_X1 U56 ( .A1(B[9]), .A2(A[9]), .ZN(n16) );
endmodule


module warp_generator_SHMEM_ADDR_SIZE14_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [3:0] A;
  input [13:0] B;
  output [17:0] PRODUCT;
  input TC;
  wire   \ab[3><13] , \ab[3><12] , \ab[3><11] , \ab[3><10] , \ab[3><9] ,
         \ab[3><8] , \ab[3><7] , \ab[3><6] , \ab[3><5] , \ab[3><4] ,
         \ab[3><3] , \ab[3><2] , \ab[3><1] , \ab[3><0] , \ab[2><13] ,
         \ab[2><12] , \ab[2><11] , \ab[2><10] , \ab[2><9] , \ab[2><8] ,
         \ab[2><7] , \ab[2><6] , \ab[2><5] , \ab[2><4] , \ab[2><3] ,
         \ab[2><2] , \ab[2><1] , \ab[2><0] , \ab[1><13] , \ab[1><12] ,
         \ab[1><11] , \ab[1><10] , \ab[1><9] , \ab[1><8] , \ab[1><7] ,
         \ab[1><6] , \ab[1><5] , \ab[1><4] , \ab[1><3] , \ab[1><2] ,
         \ab[1><1] , \ab[1><0] , \ab[0><13] , \ab[0><12] , \ab[0><11] ,
         \ab[0><10] , \ab[0><9] , \ab[0><8] , \ab[0><7] , \ab[0><6] ,
         \ab[0><5] , \ab[0><4] , \ab[0><3] , \ab[0><2] , \ab[0><1] ,
         \CARRYB[3><12] , \CARRYB[3><11] , \CARRYB[3><10] , \CARRYB[3><9] ,
         \CARRYB[3><8] , \CARRYB[3><7] , \CARRYB[3><6] , \CARRYB[3><5] ,
         \CARRYB[3><4] , \CARRYB[3><3] , \CARRYB[3><2] , \CARRYB[3><1] ,
         \CARRYB[3><0] , \CARRYB[2><12] , \CARRYB[2><11] , \CARRYB[2><10] ,
         \CARRYB[2><9] , \CARRYB[2><8] , \CARRYB[2><7] , \CARRYB[2><6] ,
         \CARRYB[2><5] , \CARRYB[2><4] , \CARRYB[2><3] , \CARRYB[2><2] ,
         \CARRYB[2><1] , \CARRYB[2><0] , \SUMB[3><12] , \SUMB[3><11] ,
         \SUMB[3><10] , \SUMB[3><9] , \SUMB[3><8] , \SUMB[3><7] , \SUMB[3><6] ,
         \SUMB[3><5] , \SUMB[3><4] , \SUMB[3><3] , \SUMB[3><2] , \SUMB[3><1] ,
         \SUMB[3><0] , \SUMB[2><12] , \SUMB[2><11] , \SUMB[2><10] ,
         \SUMB[2><9] , \SUMB[2><8] , \SUMB[2><7] , \SUMB[2><6] , \SUMB[2><5] ,
         \SUMB[2><4] , \SUMB[2><3] , \SUMB[2><2] , \SUMB[2><1] , \A1[0] , n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;

  FA_X1 S4_0 ( .A(\ab[3><0] ), .B(\CARRYB[2><0] ), .CI(\SUMB[2><1] ), .CO(
        \CARRYB[3><0] ), .S(\SUMB[3><0] ) );
  FA_X1 S4_1 ( .A(\ab[3><1] ), .B(\CARRYB[2><1] ), .CI(\SUMB[2><2] ), .CO(
        \CARRYB[3><1] ), .S(\SUMB[3><1] ) );
  FA_X1 S4_2 ( .A(\ab[3><2] ), .B(\CARRYB[2><2] ), .CI(\SUMB[2><3] ), .CO(
        \CARRYB[3><2] ), .S(\SUMB[3><2] ) );
  FA_X1 S4_3 ( .A(\ab[3><3] ), .B(\CARRYB[2><3] ), .CI(\SUMB[2><4] ), .CO(
        \CARRYB[3><3] ), .S(\SUMB[3><3] ) );
  FA_X1 S4_4 ( .A(\ab[3><4] ), .B(\CARRYB[2><4] ), .CI(\SUMB[2><5] ), .CO(
        \CARRYB[3><4] ), .S(\SUMB[3><4] ) );
  FA_X1 S4_5 ( .A(\ab[3><5] ), .B(\CARRYB[2><5] ), .CI(\SUMB[2><6] ), .CO(
        \CARRYB[3><5] ), .S(\SUMB[3><5] ) );
  FA_X1 S4_6 ( .A(\ab[3><6] ), .B(\CARRYB[2><6] ), .CI(\SUMB[2><7] ), .CO(
        \CARRYB[3><6] ), .S(\SUMB[3><6] ) );
  FA_X1 S4_7 ( .A(\ab[3><7] ), .B(\CARRYB[2><7] ), .CI(\SUMB[2><8] ), .CO(
        \CARRYB[3><7] ), .S(\SUMB[3><7] ) );
  FA_X1 S4_8 ( .A(\ab[3><8] ), .B(\CARRYB[2><8] ), .CI(\SUMB[2><9] ), .CO(
        \CARRYB[3><8] ), .S(\SUMB[3><8] ) );
  FA_X1 S4_9 ( .A(\ab[3><9] ), .B(\CARRYB[2><9] ), .CI(\SUMB[2><10] ), .CO(
        \CARRYB[3><9] ), .S(\SUMB[3><9] ) );
  FA_X1 S4_10 ( .A(\ab[3><10] ), .B(\CARRYB[2><10] ), .CI(\SUMB[2><11] ), .CO(
        \CARRYB[3><10] ), .S(\SUMB[3><10] ) );
  FA_X1 S4_11 ( .A(\ab[3><11] ), .B(\CARRYB[2><11] ), .CI(\SUMB[2><12] ), .CO(
        \CARRYB[3><11] ), .S(\SUMB[3><11] ) );
  FA_X1 S5_12 ( .A(\ab[3><12] ), .B(\CARRYB[2><12] ), .CI(\ab[2><13] ), .CO(
        \CARRYB[3><12] ), .S(\SUMB[3><12] ) );
  FA_X1 S1_2_0 ( .A(\ab[2><0] ), .B(n20), .CI(n34), .CO(\CARRYB[2><0] ), .S(
        \A1[0] ) );
  FA_X1 S2_2_1 ( .A(\ab[2><1] ), .B(n19), .CI(n33), .CO(\CARRYB[2><1] ), .S(
        \SUMB[2><1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2><2] ), .B(n18), .CI(n32), .CO(\CARRYB[2><2] ), .S(
        \SUMB[2><2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2><3] ), .B(n17), .CI(n31), .CO(\CARRYB[2><3] ), .S(
        \SUMB[2><3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2><4] ), .B(n16), .CI(n30), .CO(\CARRYB[2><4] ), .S(
        \SUMB[2><4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2><5] ), .B(n15), .CI(n29), .CO(\CARRYB[2><5] ), .S(
        \SUMB[2><5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2><6] ), .B(n14), .CI(n28), .CO(\CARRYB[2><6] ), .S(
        \SUMB[2><6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2><7] ), .B(n13), .CI(n27), .CO(\CARRYB[2><7] ), .S(
        \SUMB[2><7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2><8] ), .B(n12), .CI(n26), .CO(\CARRYB[2><8] ), .S(
        \SUMB[2><8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2><9] ), .B(n11), .CI(n25), .CO(\CARRYB[2><9] ), .S(
        \SUMB[2><9] ) );
  FA_X1 S2_2_10 ( .A(\ab[2><10] ), .B(n10), .CI(n24), .CO(\CARRYB[2><10] ), 
        .S(\SUMB[2><10] ) );
  FA_X1 S2_2_11 ( .A(\ab[2><11] ), .B(n9), .CI(n23), .CO(\CARRYB[2><11] ), .S(
        \SUMB[2><11] ) );
  FA_X1 S3_2_12 ( .A(\ab[2><12] ), .B(n37), .CI(\ab[1><13] ), .CO(
        \CARRYB[2><12] ), .S(\SUMB[2><12] ) );
  warp_generator_SHMEM_ADDR_SIZE14_DW01_add_1 FS_1 ( .A({1'b0, n2, n4, n5, n21, 
        n53, n48, n52, n47, n40, n46, n39, n38, n36, \SUMB[3><0] , \A1[0] }), 
        .B({n3, n7, n6, n8, n35, n50, n45, n49, n44, n51, n43, n42, n41, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, PRODUCT[13:2]}) );
  XOR2_X1 U2 ( .A(\CARRYB[3><12] ), .B(\ab[3><13] ), .Z(n2) );
  AND2_X1 U3 ( .A1(\CARRYB[3><12] ), .A2(\ab[3><13] ), .ZN(n3) );
  XOR2_X1 U4 ( .A(\CARRYB[3><11] ), .B(\SUMB[3><12] ), .Z(n4) );
  XOR2_X1 U5 ( .A(\CARRYB[3><10] ), .B(\SUMB[3><11] ), .Z(n5) );
  AND2_X1 U6 ( .A1(\CARRYB[3><10] ), .A2(\SUMB[3><11] ), .ZN(n6) );
  AND2_X1 U7 ( .A1(\CARRYB[3><11] ), .A2(\SUMB[3><12] ), .ZN(n7) );
  AND2_X1 U8 ( .A1(\CARRYB[3><9] ), .A2(\SUMB[3><10] ), .ZN(n8) );
  AND2_X1 U9 ( .A1(\ab[0><12] ), .A2(\ab[1><11] ), .ZN(n9) );
  AND2_X1 U10 ( .A1(\ab[0><11] ), .A2(\ab[1><10] ), .ZN(n10) );
  AND2_X1 U11 ( .A1(\ab[0><10] ), .A2(\ab[1><9] ), .ZN(n11) );
  AND2_X1 U12 ( .A1(\ab[0><9] ), .A2(\ab[1><8] ), .ZN(n12) );
  AND2_X1 U13 ( .A1(\ab[0><8] ), .A2(\ab[1><7] ), .ZN(n13) );
  AND2_X1 U14 ( .A1(\ab[0><7] ), .A2(\ab[1><6] ), .ZN(n14) );
  AND2_X1 U15 ( .A1(\ab[0><6] ), .A2(\ab[1><5] ), .ZN(n15) );
  AND2_X1 U16 ( .A1(\ab[0><5] ), .A2(\ab[1><4] ), .ZN(n16) );
  AND2_X1 U17 ( .A1(\ab[0><4] ), .A2(\ab[1><3] ), .ZN(n17) );
  AND2_X1 U18 ( .A1(\ab[0><3] ), .A2(\ab[1><2] ), .ZN(n18) );
  AND2_X1 U19 ( .A1(\ab[0><2] ), .A2(\ab[1><1] ), .ZN(n19) );
  AND2_X1 U20 ( .A1(\ab[0><1] ), .A2(\ab[1><0] ), .ZN(n20) );
  XOR2_X1 U21 ( .A(\CARRYB[3><9] ), .B(\SUMB[3><10] ), .Z(n21) );
  XOR2_X1 U22 ( .A(\ab[1><0] ), .B(\ab[0><1] ), .Z(PRODUCT[1]) );
  XOR2_X1 U23 ( .A(\ab[1><12] ), .B(\ab[0><13] ), .Z(n23) );
  XOR2_X1 U24 ( .A(\ab[1><11] ), .B(\ab[0><12] ), .Z(n24) );
  XOR2_X1 U25 ( .A(\ab[1><10] ), .B(\ab[0><11] ), .Z(n25) );
  XOR2_X1 U26 ( .A(\ab[1><9] ), .B(\ab[0><10] ), .Z(n26) );
  XOR2_X1 U27 ( .A(\ab[1><8] ), .B(\ab[0><9] ), .Z(n27) );
  XOR2_X1 U28 ( .A(\ab[1><7] ), .B(\ab[0><8] ), .Z(n28) );
  XOR2_X1 U29 ( .A(\ab[1><6] ), .B(\ab[0><7] ), .Z(n29) );
  XOR2_X1 U30 ( .A(\ab[1><5] ), .B(\ab[0><6] ), .Z(n30) );
  XOR2_X1 U31 ( .A(\ab[1><4] ), .B(\ab[0><5] ), .Z(n31) );
  XOR2_X1 U32 ( .A(\ab[1><3] ), .B(\ab[0><4] ), .Z(n32) );
  XOR2_X1 U33 ( .A(\ab[1><2] ), .B(\ab[0><3] ), .Z(n33) );
  XOR2_X1 U34 ( .A(\ab[1><1] ), .B(\ab[0><2] ), .Z(n34) );
  AND2_X1 U35 ( .A1(\CARRYB[3><8] ), .A2(\SUMB[3><9] ), .ZN(n35) );
  XOR2_X1 U36 ( .A(\CARRYB[3><0] ), .B(\SUMB[3><1] ), .Z(n36) );
  AND2_X1 U37 ( .A1(\ab[0><13] ), .A2(\ab[1><12] ), .ZN(n37) );
  XOR2_X1 U38 ( .A(\CARRYB[3><1] ), .B(\SUMB[3><2] ), .Z(n38) );
  XOR2_X1 U39 ( .A(\CARRYB[3><2] ), .B(\SUMB[3><3] ), .Z(n39) );
  XOR2_X1 U40 ( .A(\CARRYB[3><4] ), .B(\SUMB[3><5] ), .Z(n40) );
  AND2_X1 U41 ( .A1(\CARRYB[3><0] ), .A2(\SUMB[3><1] ), .ZN(n41) );
  AND2_X1 U42 ( .A1(\CARRYB[3><1] ), .A2(\SUMB[3><2] ), .ZN(n42) );
  AND2_X1 U43 ( .A1(\CARRYB[3><2] ), .A2(\SUMB[3><3] ), .ZN(n43) );
  AND2_X1 U44 ( .A1(\CARRYB[3><4] ), .A2(\SUMB[3><5] ), .ZN(n44) );
  AND2_X1 U45 ( .A1(\CARRYB[3><6] ), .A2(\SUMB[3><7] ), .ZN(n45) );
  XOR2_X1 U46 ( .A(\CARRYB[3><3] ), .B(\SUMB[3><4] ), .Z(n46) );
  XOR2_X1 U47 ( .A(\CARRYB[3><5] ), .B(\SUMB[3><6] ), .Z(n47) );
  XOR2_X1 U48 ( .A(\CARRYB[3><7] ), .B(\SUMB[3><8] ), .Z(n48) );
  AND2_X1 U49 ( .A1(\CARRYB[3><5] ), .A2(\SUMB[3><6] ), .ZN(n49) );
  AND2_X1 U50 ( .A1(\CARRYB[3><7] ), .A2(\SUMB[3><8] ), .ZN(n50) );
  AND2_X1 U51 ( .A1(\CARRYB[3><3] ), .A2(\SUMB[3><4] ), .ZN(n51) );
  XOR2_X1 U52 ( .A(\CARRYB[3><6] ), .B(\SUMB[3><7] ), .Z(n52) );
  XOR2_X1 U53 ( .A(\CARRYB[3><8] ), .B(\SUMB[3><9] ), .Z(n53) );
  INV_X1 U54 ( .A(A[1]), .ZN(n55) );
  INV_X1 U55 ( .A(A[3]), .ZN(n57) );
  INV_X1 U56 ( .A(A[0]), .ZN(n54) );
  INV_X1 U57 ( .A(A[2]), .ZN(n56) );
  INV_X1 U58 ( .A(B[1]), .ZN(n70) );
  INV_X1 U59 ( .A(B[0]), .ZN(n71) );
  INV_X1 U60 ( .A(B[2]), .ZN(n69) );
  INV_X1 U61 ( .A(B[3]), .ZN(n68) );
  INV_X1 U62 ( .A(B[6]), .ZN(n65) );
  INV_X1 U63 ( .A(B[4]), .ZN(n67) );
  INV_X1 U64 ( .A(B[5]), .ZN(n66) );
  INV_X1 U65 ( .A(B[8]), .ZN(n63) );
  INV_X1 U66 ( .A(B[7]), .ZN(n64) );
  INV_X1 U67 ( .A(B[10]), .ZN(n61) );
  INV_X1 U68 ( .A(B[9]), .ZN(n62) );
  INV_X1 U69 ( .A(B[11]), .ZN(n60) );
  INV_X1 U70 ( .A(B[12]), .ZN(n59) );
  INV_X1 U71 ( .A(B[13]), .ZN(n58) );
  NOR2_X1 U73 ( .A1(n57), .A2(n62), .ZN(\ab[3><9] ) );
  NOR2_X1 U74 ( .A1(n57), .A2(n63), .ZN(\ab[3><8] ) );
  NOR2_X1 U75 ( .A1(n57), .A2(n64), .ZN(\ab[3><7] ) );
  NOR2_X1 U76 ( .A1(n57), .A2(n65), .ZN(\ab[3><6] ) );
  NOR2_X1 U77 ( .A1(n57), .A2(n66), .ZN(\ab[3><5] ) );
  NOR2_X1 U78 ( .A1(n57), .A2(n67), .ZN(\ab[3><4] ) );
  NOR2_X1 U79 ( .A1(n57), .A2(n68), .ZN(\ab[3><3] ) );
  NOR2_X1 U80 ( .A1(n57), .A2(n69), .ZN(\ab[3><2] ) );
  NOR2_X1 U81 ( .A1(n57), .A2(n70), .ZN(\ab[3><1] ) );
  NOR2_X1 U82 ( .A1(n57), .A2(n58), .ZN(\ab[3><13] ) );
  NOR2_X1 U83 ( .A1(n57), .A2(n59), .ZN(\ab[3><12] ) );
  NOR2_X1 U84 ( .A1(n57), .A2(n60), .ZN(\ab[3><11] ) );
  NOR2_X1 U85 ( .A1(n57), .A2(n61), .ZN(\ab[3><10] ) );
  NOR2_X1 U86 ( .A1(n57), .A2(n71), .ZN(\ab[3><0] ) );
  NOR2_X1 U87 ( .A1(n62), .A2(n56), .ZN(\ab[2><9] ) );
  NOR2_X1 U88 ( .A1(n63), .A2(n56), .ZN(\ab[2><8] ) );
  NOR2_X1 U89 ( .A1(n64), .A2(n56), .ZN(\ab[2><7] ) );
  NOR2_X1 U90 ( .A1(n65), .A2(n56), .ZN(\ab[2><6] ) );
  NOR2_X1 U91 ( .A1(n66), .A2(n56), .ZN(\ab[2><5] ) );
  NOR2_X1 U92 ( .A1(n67), .A2(n56), .ZN(\ab[2><4] ) );
  NOR2_X1 U93 ( .A1(n68), .A2(n56), .ZN(\ab[2><3] ) );
  NOR2_X1 U94 ( .A1(n69), .A2(n56), .ZN(\ab[2><2] ) );
  NOR2_X1 U95 ( .A1(n70), .A2(n56), .ZN(\ab[2><1] ) );
  NOR2_X1 U96 ( .A1(n58), .A2(n56), .ZN(\ab[2><13] ) );
  NOR2_X1 U97 ( .A1(n59), .A2(n56), .ZN(\ab[2><12] ) );
  NOR2_X1 U98 ( .A1(n60), .A2(n56), .ZN(\ab[2><11] ) );
  NOR2_X1 U99 ( .A1(n61), .A2(n56), .ZN(\ab[2><10] ) );
  NOR2_X1 U100 ( .A1(n71), .A2(n56), .ZN(\ab[2><0] ) );
  NOR2_X1 U101 ( .A1(n62), .A2(n55), .ZN(\ab[1><9] ) );
  NOR2_X1 U102 ( .A1(n63), .A2(n55), .ZN(\ab[1><8] ) );
  NOR2_X1 U103 ( .A1(n64), .A2(n55), .ZN(\ab[1><7] ) );
  NOR2_X1 U104 ( .A1(n65), .A2(n55), .ZN(\ab[1><6] ) );
  NOR2_X1 U105 ( .A1(n66), .A2(n55), .ZN(\ab[1><5] ) );
  NOR2_X1 U106 ( .A1(n67), .A2(n55), .ZN(\ab[1><4] ) );
  NOR2_X1 U107 ( .A1(n68), .A2(n55), .ZN(\ab[1><3] ) );
  NOR2_X1 U108 ( .A1(n69), .A2(n55), .ZN(\ab[1><2] ) );
  NOR2_X1 U109 ( .A1(n70), .A2(n55), .ZN(\ab[1><1] ) );
  NOR2_X1 U110 ( .A1(n58), .A2(n55), .ZN(\ab[1><13] ) );
  NOR2_X1 U111 ( .A1(n59), .A2(n55), .ZN(\ab[1><12] ) );
  NOR2_X1 U112 ( .A1(n60), .A2(n55), .ZN(\ab[1><11] ) );
  NOR2_X1 U113 ( .A1(n61), .A2(n55), .ZN(\ab[1><10] ) );
  NOR2_X1 U114 ( .A1(n71), .A2(n55), .ZN(\ab[1><0] ) );
  NOR2_X1 U115 ( .A1(n62), .A2(n54), .ZN(\ab[0><9] ) );
  NOR2_X1 U116 ( .A1(n63), .A2(n54), .ZN(\ab[0><8] ) );
  NOR2_X1 U117 ( .A1(n64), .A2(n54), .ZN(\ab[0><7] ) );
  NOR2_X1 U118 ( .A1(n65), .A2(n54), .ZN(\ab[0><6] ) );
  NOR2_X1 U119 ( .A1(n66), .A2(n54), .ZN(\ab[0><5] ) );
  NOR2_X1 U120 ( .A1(n67), .A2(n54), .ZN(\ab[0><4] ) );
  NOR2_X1 U121 ( .A1(n68), .A2(n54), .ZN(\ab[0><3] ) );
  NOR2_X1 U122 ( .A1(n69), .A2(n54), .ZN(\ab[0><2] ) );
  NOR2_X1 U123 ( .A1(n70), .A2(n54), .ZN(\ab[0><1] ) );
  NOR2_X1 U124 ( .A1(n58), .A2(n54), .ZN(\ab[0><13] ) );
  NOR2_X1 U125 ( .A1(n59), .A2(n54), .ZN(\ab[0><12] ) );
  NOR2_X1 U126 ( .A1(n60), .A2(n54), .ZN(\ab[0><11] ) );
  NOR2_X1 U127 ( .A1(n61), .A2(n54), .ZN(\ab[0><10] ) );
  NOR2_X1 U128 ( .A1(n71), .A2(n54), .ZN(PRODUCT[0]) );
endmodule



module warp_generator_SHMEM_ADDR_SIZE14_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [13:1] carry;

  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .S(SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(n2) );
endmodule



module warp_generator ( clk_in, host_reset, en, 
        num_blocks_in, warps_per_block_in, shmem_base_addr_in, shmem_size_in, 
        gprs_size_in, warp_pool_addr_out, warp_pool_wr_en_out, 
        warp_pool_wr_data_out, warp_state_addr_out, warp_state_wr_en_out, 
        warp_state_wr_data_out, .fence_regs_cta_id_out({
        \fence_regs_cta_id_out[31><3] , \fence_regs_cta_id_out[31><2] , 
        \fence_regs_cta_id_out[31><1] , \fence_regs_cta_id_out[31><0] , 
        \fence_regs_cta_id_out[30><3] , \fence_regs_cta_id_out[30><2] , 
        \fence_regs_cta_id_out[30><1] , \fence_regs_cta_id_out[30><0] , 
        \fence_regs_cta_id_out[29><3] , \fence_regs_cta_id_out[29><2] , 
        \fence_regs_cta_id_out[29><1] , \fence_regs_cta_id_out[29><0] , 
        \fence_regs_cta_id_out[28><3] , \fence_regs_cta_id_out[28><2] , 
        \fence_regs_cta_id_out[28><1] , \fence_regs_cta_id_out[28><0] , 
        \fence_regs_cta_id_out[27><3] , \fence_regs_cta_id_out[27><2] , 
        \fence_regs_cta_id_out[27><1] , \fence_regs_cta_id_out[27><0] , 
        \fence_regs_cta_id_out[26><3] , \fence_regs_cta_id_out[26><2] , 
        \fence_regs_cta_id_out[26><1] , \fence_regs_cta_id_out[26><0] , 
        \fence_regs_cta_id_out[25><3] , \fence_regs_cta_id_out[25><2] , 
        \fence_regs_cta_id_out[25><1] , \fence_regs_cta_id_out[25><0] , 
        \fence_regs_cta_id_out[24><3] , \fence_regs_cta_id_out[24><2] , 
        \fence_regs_cta_id_out[24><1] , \fence_regs_cta_id_out[24><0] , 
        \fence_regs_cta_id_out[23><3] , \fence_regs_cta_id_out[23><2] , 
        \fence_regs_cta_id_out[23><1] , \fence_regs_cta_id_out[23><0] , 
        \fence_regs_cta_id_out[22><3] , \fence_regs_cta_id_out[22><2] , 
        \fence_regs_cta_id_out[22><1] , \fence_regs_cta_id_out[22><0] , 
        \fence_regs_cta_id_out[21><3] , \fence_regs_cta_id_out[21><2] , 
        \fence_regs_cta_id_out[21><1] , \fence_regs_cta_id_out[21><0] , 
        \fence_regs_cta_id_out[20><3] , \fence_regs_cta_id_out[20><2] , 
        \fence_regs_cta_id_out[20><1] , \fence_regs_cta_id_out[20><0] , 
        \fence_regs_cta_id_out[19><3] , \fence_regs_cta_id_out[19><2] , 
        \fence_regs_cta_id_out[19><1] , \fence_regs_cta_id_out[19><0] , 
        \fence_regs_cta_id_out[18><3] , \fence_regs_cta_id_out[18><2] , 
        \fence_regs_cta_id_out[18><1] , \fence_regs_cta_id_out[18><0] , 
        \fence_regs_cta_id_out[17><3] , \fence_regs_cta_id_out[17><2] , 
        \fence_regs_cta_id_out[17><1] , \fence_regs_cta_id_out[17><0] , 
        \fence_regs_cta_id_out[16><3] , \fence_regs_cta_id_out[16><2] , 
        \fence_regs_cta_id_out[16><1] , \fence_regs_cta_id_out[16><0] , 
        \fence_regs_cta_id_out[15><3] , \fence_regs_cta_id_out[15><2] , 
        \fence_regs_cta_id_out[15><1] , \fence_regs_cta_id_out[15><0] , 
        \fence_regs_cta_id_out[14><3] , \fence_regs_cta_id_out[14><2] , 
        \fence_regs_cta_id_out[14><1] , \fence_regs_cta_id_out[14><0] , 
        \fence_regs_cta_id_out[13><3] , \fence_regs_cta_id_out[13><2] , 
        \fence_regs_cta_id_out[13><1] , \fence_regs_cta_id_out[13><0] , 
        \fence_regs_cta_id_out[12><3] , \fence_regs_cta_id_out[12><2] , 
        \fence_regs_cta_id_out[12><1] , \fence_regs_cta_id_out[12><0] , 
        \fence_regs_cta_id_out[11><3] , \fence_regs_cta_id_out[11><2] , 
        \fence_regs_cta_id_out[11><1] , \fence_regs_cta_id_out[11><0] , 
        \fence_regs_cta_id_out[10><3] , \fence_regs_cta_id_out[10><2] , 
        \fence_regs_cta_id_out[10><1] , \fence_regs_cta_id_out[10><0] , 
        \fence_regs_cta_id_out[9><3] , \fence_regs_cta_id_out[9><2] , 
        \fence_regs_cta_id_out[9><1] , \fence_regs_cta_id_out[9><0] , 
        \fence_regs_cta_id_out[8><3] , \fence_regs_cta_id_out[8><2] , 
        \fence_regs_cta_id_out[8><1] , \fence_regs_cta_id_out[8><0] , 
        \fence_regs_cta_id_out[7><3] , \fence_regs_cta_id_out[7><2] , 
        \fence_regs_cta_id_out[7><1] , \fence_regs_cta_id_out[7><0] , 
        \fence_regs_cta_id_out[6><3] , \fence_regs_cta_id_out[6><2] , 
        \fence_regs_cta_id_out[6><1] , \fence_regs_cta_id_out[6><0] , 
        \fence_regs_cta_id_out[5><3] , \fence_regs_cta_id_out[5><2] , 
        \fence_regs_cta_id_out[5><1] , \fence_regs_cta_id_out[5><0] , 
        \fence_regs_cta_id_out[4><3] , \fence_regs_cta_id_out[4><2] , 
        \fence_regs_cta_id_out[4><1] , \fence_regs_cta_id_out[4><0] , 
        \fence_regs_cta_id_out[3><3] , \fence_regs_cta_id_out[3><2] , 
        \fence_regs_cta_id_out[3><1] , \fence_regs_cta_id_out[3><0] , 
        \fence_regs_cta_id_out[2><3] , \fence_regs_cta_id_out[2><2] , 
        \fence_regs_cta_id_out[2><1] , \fence_regs_cta_id_out[2><0] , 
        \fence_regs_cta_id_out[1><3] , \fence_regs_cta_id_out[1><2] , 
        \fence_regs_cta_id_out[1><1] , \fence_regs_cta_id_out[1><0] , 
        \fence_regs_cta_id_out[0><3] , \fence_regs_cta_id_out[0><2] , 
        \fence_regs_cta_id_out[0><1] , \fence_regs_cta_id_out[0><0] }), 
        fence_regs_cta_id_ld, fence_regs_fence_en_out, fence_regs_fence_en_ld, 
        num_warps_out, warp_gen_done );
  input [3:0] num_blocks_in;
  input [5:0] warps_per_block_in;
  input [31:0] shmem_base_addr_in;
  input [31:0] shmem_size_in;
  input [8:0] gprs_size_in;
  output [4:0] warp_pool_addr_out;
  output [127:0] warp_pool_wr_data_out;
  output [4:0] warp_state_addr_out;
  output [1:0] warp_state_wr_data_out;
  output [31:0] fence_regs_cta_id_ld;
  output [31:0] fence_regs_fence_en_out;
  output [31:0] fence_regs_fence_en_ld;
  output [4:0] num_warps_out;
  input clk_in, host_reset, en;
  output warp_pool_wr_en_out, warp_state_wr_en_out,
         \fence_regs_cta_id_out[31><3] , \fence_regs_cta_id_out[31><2] ,
         \fence_regs_cta_id_out[31><1] , \fence_regs_cta_id_out[31><0] ,
         \fence_regs_cta_id_out[30><3] , \fence_regs_cta_id_out[30><2] ,
         \fence_regs_cta_id_out[30><1] , \fence_regs_cta_id_out[30><0] ,
         \fence_regs_cta_id_out[29><3] , \fence_regs_cta_id_out[29><2] ,
         \fence_regs_cta_id_out[29><1] , \fence_regs_cta_id_out[29><0] ,
         \fence_regs_cta_id_out[28><3] , \fence_regs_cta_id_out[28><2] ,
         \fence_regs_cta_id_out[28><1] , \fence_regs_cta_id_out[28><0] ,
         \fence_regs_cta_id_out[27><3] , \fence_regs_cta_id_out[27><2] ,
         \fence_regs_cta_id_out[27><1] , \fence_regs_cta_id_out[27><0] ,
         \fence_regs_cta_id_out[26><3] , \fence_regs_cta_id_out[26><2] ,
         \fence_regs_cta_id_out[26><1] , \fence_regs_cta_id_out[26><0] ,
         \fence_regs_cta_id_out[25><3] , \fence_regs_cta_id_out[25><2] ,
         \fence_regs_cta_id_out[25><1] , \fence_regs_cta_id_out[25><0] ,
         \fence_regs_cta_id_out[24><3] , \fence_regs_cta_id_out[24><2] ,
         \fence_regs_cta_id_out[24><1] , \fence_regs_cta_id_out[24><0] ,
         \fence_regs_cta_id_out[23><3] , \fence_regs_cta_id_out[23><2] ,
         \fence_regs_cta_id_out[23><1] , \fence_regs_cta_id_out[23><0] ,
         \fence_regs_cta_id_out[22><3] , \fence_regs_cta_id_out[22><2] ,
         \fence_regs_cta_id_out[22><1] , \fence_regs_cta_id_out[22><0] ,
         \fence_regs_cta_id_out[21><3] , \fence_regs_cta_id_out[21><2] ,
         \fence_regs_cta_id_out[21><1] , \fence_regs_cta_id_out[21><0] ,
         \fence_regs_cta_id_out[20><3] , \fence_regs_cta_id_out[20><2] ,
         \fence_regs_cta_id_out[20><1] , \fence_regs_cta_id_out[20><0] ,
         \fence_regs_cta_id_out[19><3] , \fence_regs_cta_id_out[19><2] ,
         \fence_regs_cta_id_out[19><1] , \fence_regs_cta_id_out[19><0] ,
         \fence_regs_cta_id_out[18><3] , \fence_regs_cta_id_out[18><2] ,
         \fence_regs_cta_id_out[18><1] , \fence_regs_cta_id_out[18><0] ,
         \fence_regs_cta_id_out[17><3] , \fence_regs_cta_id_out[17><2] ,
         \fence_regs_cta_id_out[17><1] , \fence_regs_cta_id_out[17><0] ,
         \fence_regs_cta_id_out[16><3] , \fence_regs_cta_id_out[16><2] ,
         \fence_regs_cta_id_out[16><1] , \fence_regs_cta_id_out[16><0] ,
         \fence_regs_cta_id_out[15><3] , \fence_regs_cta_id_out[15><2] ,
         \fence_regs_cta_id_out[15><1] , \fence_regs_cta_id_out[15><0] ,
         \fence_regs_cta_id_out[14><3] , \fence_regs_cta_id_out[14><2] ,
         \fence_regs_cta_id_out[14><1] , \fence_regs_cta_id_out[14><0] ,
         \fence_regs_cta_id_out[13><3] , \fence_regs_cta_id_out[13><2] ,
         \fence_regs_cta_id_out[13><1] , \fence_regs_cta_id_out[13><0] ,
         \fence_regs_cta_id_out[12><3] , \fence_regs_cta_id_out[12><2] ,
         \fence_regs_cta_id_out[12><1] , \fence_regs_cta_id_out[12><0] ,
         \fence_regs_cta_id_out[11><3] , \fence_regs_cta_id_out[11><2] ,
         \fence_regs_cta_id_out[11><1] , \fence_regs_cta_id_out[11><0] ,
         \fence_regs_cta_id_out[10><3] , \fence_regs_cta_id_out[10><2] ,
         \fence_regs_cta_id_out[10><1] , \fence_regs_cta_id_out[10><0] ,
         \fence_regs_cta_id_out[9><3] , \fence_regs_cta_id_out[9><2] ,
         \fence_regs_cta_id_out[9><1] , \fence_regs_cta_id_out[9><0] ,
         \fence_regs_cta_id_out[8><3] , \fence_regs_cta_id_out[8><2] ,
         \fence_regs_cta_id_out[8><1] , \fence_regs_cta_id_out[8><0] ,
         \fence_regs_cta_id_out[7><3] , \fence_regs_cta_id_out[7><2] ,
         \fence_regs_cta_id_out[7><1] , \fence_regs_cta_id_out[7><0] ,
         \fence_regs_cta_id_out[6><3] , \fence_regs_cta_id_out[6><2] ,
         \fence_regs_cta_id_out[6><1] , \fence_regs_cta_id_out[6><0] ,
         \fence_regs_cta_id_out[5><3] , \fence_regs_cta_id_out[5><2] ,
         \fence_regs_cta_id_out[5><1] , \fence_regs_cta_id_out[5><0] ,
         \fence_regs_cta_id_out[4><3] , \fence_regs_cta_id_out[4><2] ,
         \fence_regs_cta_id_out[4><1] , \fence_regs_cta_id_out[4><0] ,
         \fence_regs_cta_id_out[3><3] , \fence_regs_cta_id_out[3><2] ,
         \fence_regs_cta_id_out[3><1] , \fence_regs_cta_id_out[3><0] ,
         \fence_regs_cta_id_out[2><3] , \fence_regs_cta_id_out[2><2] ,
         \fence_regs_cta_id_out[2><1] , \fence_regs_cta_id_out[2><0] ,
         \fence_regs_cta_id_out[1><3] , \fence_regs_cta_id_out[1><2] ,
         \fence_regs_cta_id_out[1><1] , \fence_regs_cta_id_out[1><0] ,
         \fence_regs_cta_id_out[0><3] , \fence_regs_cta_id_out[0><2] ,
         \fence_regs_cta_id_out[0><1] , \fence_regs_cta_id_out[0><0] ,
         warp_gen_done;
  wire   warp_id_calc_en_i, N62, N78, N79, N80, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N254, N255, N256, N257, N863, N864, N865, N866,
         N867, N868, N869, N870, N871, N872, N873, N874, N875, N876, N877,
         N878, N879, N880, N881, N882, N883, N884, N885, N886, N887, N888,
         N889, N890, N891, N892, N893, N894, n40, n41, n42, n43, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n141, n142, n143, n145,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, N77, N76, N75, N74, N73, N72, N71, N70, N69, N68, N67,
         N66, N65, N64, \add_155/carry[4] , \add_155/carry[3] ,
         \add_155/carry[2] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n144, n146, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n272, n273,
         n274, n275, n276, n277, n278, n279, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876;
  wire   [3:0] block_num_cnt;
  wire   [11:0] warps_per_block_cnt;
  wire   [3:0] block_num_i;
  wire   [4:0] warp_num_i;
  wire   [2:0] warp_generator_state_machine;
  wire   [13:0] shmem_addr_i;
  wire   [4:0] warp_id_o;
  wire   [4:0] warp_id_addr;
  wire   [8:0] gprs_base_addr_o;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign warp_pool_wr_data_out[127] = 1'b0;
  assign warp_pool_wr_data_out[126] = 1'b0;
  assign warp_pool_wr_data_out[125] = 1'b0;
  assign warp_pool_wr_data_out[124] = 1'b0;
  assign warp_pool_wr_data_out[96] = 1'b0;
  assign warp_pool_wr_data_out[95] = 1'b0;
  assign warp_pool_wr_data_out[94] = 1'b0;
  assign warp_pool_wr_data_out[93] = 1'b0;
  assign warp_pool_wr_data_out[92] = 1'b0;
  assign warp_pool_wr_data_out[91] = 1'b0;
  assign warp_pool_wr_data_out[90] = 1'b0;
  assign warp_pool_wr_data_out[89] = 1'b0;
  assign warp_pool_wr_data_out[88] = 1'b0;
  assign warp_pool_wr_data_out[87] = 1'b0;
  assign warp_pool_wr_data_out[86] = 1'b0;
  assign warp_pool_wr_data_out[85] = 1'b0;
  assign warp_pool_wr_data_out[84] = 1'b0;
  assign warp_pool_wr_data_out[83] = 1'b0;
  assign warp_pool_wr_data_out[82] = 1'b0;
  assign warp_pool_wr_data_out[81] = 1'b0;
  assign warp_pool_wr_data_out[80] = 1'b0;
  assign warp_pool_wr_data_out[79] = 1'b0;
  assign warp_pool_wr_data_out[78] = 1'b0;
  assign warp_pool_wr_data_out[77] = 1'b0;
  assign warp_pool_wr_data_out[76] = 1'b0;
  assign warp_pool_wr_data_out[75] = 1'b0;
  assign warp_pool_wr_data_out[74] = 1'b0;
  assign warp_pool_wr_data_out[73] = 1'b0;
  assign warp_pool_wr_data_out[72] = 1'b0;
  assign warp_pool_wr_data_out[71] = 1'b0;
  assign warp_pool_wr_data_out[70] = 1'b0;
  assign warp_pool_wr_data_out[69] = 1'b0;
  assign warp_pool_wr_data_out[68] = 1'b0;
  assign warp_pool_wr_data_out[67] = 1'b0;
  assign warp_pool_wr_data_out[66] = 1'b0;
  assign warp_pool_wr_data_out[65] = 1'b0;
  assign warp_pool_wr_data_out[64] = 1'b0;
  assign warp_state_wr_data_out[1] = 1'b0;
  assign warp_state_wr_data_out[0] = 1'b0;
  assign fence_regs_fence_en_out[31] = 1'b0;
  assign fence_regs_fence_en_out[30] = 1'b0;
  assign fence_regs_fence_en_out[29] = 1'b0;
  assign fence_regs_fence_en_out[28] = 1'b0;
  assign fence_regs_fence_en_out[27] = 1'b0;
  assign fence_regs_fence_en_out[26] = 1'b0;
  assign fence_regs_fence_en_out[25] = 1'b0;
  assign fence_regs_fence_en_out[24] = 1'b0;
  assign fence_regs_fence_en_out[23] = 1'b0;
  assign fence_regs_fence_en_out[22] = 1'b0;
  assign fence_regs_fence_en_out[21] = 1'b0;
  assign fence_regs_fence_en_out[20] = 1'b0;
  assign fence_regs_fence_en_out[19] = 1'b0;
  assign fence_regs_fence_en_out[18] = 1'b0;
  assign fence_regs_fence_en_out[17] = 1'b0;
  assign fence_regs_fence_en_out[16] = 1'b0;
  assign fence_regs_fence_en_out[15] = 1'b0;
  assign fence_regs_fence_en_out[14] = 1'b0;
  assign fence_regs_fence_en_out[13] = 1'b0;
  assign fence_regs_fence_en_out[12] = 1'b0;
  assign fence_regs_fence_en_out[11] = 1'b0;
  assign fence_regs_fence_en_out[10] = 1'b0;
  assign fence_regs_fence_en_out[9] = 1'b0;
  assign fence_regs_fence_en_out[8] = 1'b0;
  assign fence_regs_fence_en_out[7] = 1'b0;
  assign fence_regs_fence_en_out[6] = 1'b0;
  assign fence_regs_fence_en_out[5] = 1'b0;
  assign fence_regs_fence_en_out[4] = 1'b0;
  assign fence_regs_fence_en_out[3] = 1'b0;
  assign fence_regs_fence_en_out[2] = 1'b0;
  assign fence_regs_fence_en_out[1] = 1'b0;
  assign fence_regs_fence_en_out[0] = 1'b0;

  DFFR_X1 \warp_generator_state_machine_reg[0]  ( .D(n815), .CK(clk_in), .RN(
        n121), .Q(warp_generator_state_machine[0]), .QN(n202) );
  DFFR_X1 \warp_generator_state_machine_reg[1]  ( .D(n814), .CK(clk_in), .RN(
        n121), .Q(warp_generator_state_machine[1]), .QN(n201) );
  DFFR_X1 \warps_per_block_cnt_reg[11]  ( .D(n277), .CK(clk_in), .RN(n121), 
        .Q(warps_per_block_cnt[11]) );
  DFFR_X1 \warps_per_block_cnt_reg[0]  ( .D(n278), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[0]), .QN(n151) );
  DFFR_X1 \warps_per_block_cnt_reg[1]  ( .D(n279), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[1]), .QN(n150) );
  DFFR_X1 \warps_per_block_cnt_reg[2]  ( .D(n816), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[2]), .QN(n149) );
  DFFR_X1 \warps_per_block_cnt_reg[3]  ( .D(n817), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[3]), .QN(n148) );
  DFFR_X1 \warps_per_block_cnt_reg[4]  ( .D(n818), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[4]), .QN(n147) );
  DFFR_X1 \warps_per_block_cnt_reg[5]  ( .D(n819), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[5]), .QN(n2) );
  DFFR_X1 \warps_per_block_cnt_reg[6]  ( .D(n820), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[6]) );
  DFFR_X1 \warps_per_block_cnt_reg[7]  ( .D(n821), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[7]) );
  DFFR_X1 \warps_per_block_cnt_reg[8]  ( .D(n822), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[8]) );
  DFFR_X1 \warps_per_block_cnt_reg[9]  ( .D(n823), .CK(clk_in), .RN(n121), .Q(
        warps_per_block_cnt[9]) );
  DFFR_X1 \warps_per_block_cnt_reg[10]  ( .D(n824), .CK(clk_in), .RN(n121), 
        .Q(warps_per_block_cnt[10]) );
  DFFR_X1 \block_num_cnt_reg[0]  ( .D(n810), .CK(clk_in), .RN(n121), .Q(
        block_num_cnt[0]), .QN(n145) );
  DFFR_X1 \block_num_cnt_reg[1]  ( .D(n811), .CK(clk_in), .RN(n121), .Q(
        block_num_cnt[1]), .QN(n143) );
  DFFR_X1 \block_num_cnt_reg[2]  ( .D(n809), .CK(clk_in), .RN(n121), .Q(
        block_num_cnt[2]), .QN(n142) );
  DFFR_X1 \block_num_cnt_reg[3]  ( .D(n808), .CK(clk_in), .RN(n121), .Q(
        block_num_cnt[3]), .QN(n141) );
  DFFR_X1 \warp_generator_state_machine_reg[2]  ( .D(n197), .CK(clk_in), .RN(
        n122), .Q(warp_generator_state_machine[2]), .QN(n200) );
  DFFR_X1 warp_state_wr_en_out_reg ( .D(n812), .CK(clk_in), .RN(n122), .Q(
        warp_state_wr_en_out) );
  DFFR_X1 warp_pool_wr_en_out_reg ( .D(n813), .CK(clk_in), .RN(n122), .Q(
        warp_pool_wr_en_out) );
  DFFR_X1 \warp_pool_wr_data_out_reg[0]  ( .D(n733), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[0]), .QN(n116) );
  DFFR_X1 \warp_pool_wr_data_out_reg[63]  ( .D(n734), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[63]), .QN(n53) );
  DFFR_X1 \warp_pool_wr_data_out_reg[62]  ( .D(n735), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[62]), .QN(n54) );
  DFFR_X1 \warp_pool_wr_data_out_reg[61]  ( .D(n736), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[61]), .QN(n55) );
  DFFR_X1 \warp_pool_wr_data_out_reg[60]  ( .D(n737), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[60]), .QN(n56) );
  DFFR_X1 \warp_pool_wr_data_out_reg[59]  ( .D(n738), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[59]), .QN(n57) );
  DFFR_X1 \warp_pool_wr_data_out_reg[58]  ( .D(n739), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[58]), .QN(n58) );
  DFFR_X1 \warp_pool_wr_data_out_reg[57]  ( .D(n740), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[57]), .QN(n59) );
  DFFR_X1 \warp_pool_wr_data_out_reg[56]  ( .D(n741), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[56]), .QN(n60) );
  DFFR_X1 \warp_pool_wr_data_out_reg[55]  ( .D(n742), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[55]), .QN(n61) );
  DFFR_X1 \warp_pool_wr_data_out_reg[54]  ( .D(n743), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[54]), .QN(n62) );
  DFFR_X1 \warp_pool_wr_data_out_reg[53]  ( .D(n744), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[53]), .QN(n63) );
  DFFR_X1 \warp_pool_wr_data_out_reg[52]  ( .D(n745), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[52]), .QN(n64) );
  DFFR_X1 \warp_pool_wr_data_out_reg[51]  ( .D(n746), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[51]), .QN(n65) );
  DFFR_X1 \warp_pool_wr_data_out_reg[50]  ( .D(n747), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[50]), .QN(n66) );
  DFFR_X1 \warp_pool_wr_data_out_reg[49]  ( .D(n748), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[49]), .QN(n67) );
  DFFR_X1 \warp_pool_wr_data_out_reg[48]  ( .D(n749), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[48]), .QN(n68) );
  DFFR_X1 \warp_pool_wr_data_out_reg[47]  ( .D(n750), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[47]), .QN(n69) );
  DFFR_X1 \warp_pool_wr_data_out_reg[46]  ( .D(n751), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[46]), .QN(n70) );
  DFFR_X1 \warp_pool_wr_data_out_reg[45]  ( .D(n752), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[45]), .QN(n71) );
  DFFR_X1 \warp_pool_wr_data_out_reg[44]  ( .D(n753), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[44]), .QN(n72) );
  DFFR_X1 \warp_pool_wr_data_out_reg[43]  ( .D(n754), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[43]), .QN(n73) );
  DFFR_X1 \warp_pool_wr_data_out_reg[42]  ( .D(n755), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[42]), .QN(n74) );
  DFFR_X1 \warp_pool_wr_data_out_reg[41]  ( .D(n756), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[41]), .QN(n75) );
  DFFR_X1 \warp_pool_wr_data_out_reg[40]  ( .D(n757), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[40]), .QN(n76) );
  DFFR_X1 \warp_pool_wr_data_out_reg[39]  ( .D(n758), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[39]), .QN(n77) );
  DFFR_X1 \warp_pool_wr_data_out_reg[38]  ( .D(n759), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[38]), .QN(n78) );
  DFFR_X1 \warp_pool_wr_data_out_reg[37]  ( .D(n760), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[37]), .QN(n79) );
  DFFR_X1 \warp_pool_wr_data_out_reg[36]  ( .D(n761), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[36]), .QN(n80) );
  DFFR_X1 \warp_pool_wr_data_out_reg[35]  ( .D(n762), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[35]), .QN(n81) );
  DFFR_X1 \warp_pool_wr_data_out_reg[34]  ( .D(n763), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[34]), .QN(n82) );
  DFFR_X1 \warp_pool_wr_data_out_reg[33]  ( .D(n764), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[33]), .QN(n83) );
  DFFR_X1 \warp_pool_wr_data_out_reg[32]  ( .D(n765), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[32]), .QN(n84) );
  DFFR_X1 \warp_pool_wr_data_out_reg[31]  ( .D(n766), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[31]), .QN(n85) );
  DFFR_X1 \warp_pool_wr_data_out_reg[30]  ( .D(n767), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[30]), .QN(n86) );
  DFFR_X1 \warp_pool_wr_data_out_reg[29]  ( .D(n768), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[29]), .QN(n87) );
  DFFR_X1 \warp_pool_wr_data_out_reg[28]  ( .D(n769), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[28]), .QN(n88) );
  DFFR_X1 \warp_pool_wr_data_out_reg[27]  ( .D(n770), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[27]), .QN(n89) );
  DFFR_X1 \warp_pool_wr_data_out_reg[26]  ( .D(n771), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[26]), .QN(n90) );
  DFFR_X1 \warp_pool_wr_data_out_reg[25]  ( .D(n772), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[25]), .QN(n91) );
  DFFR_X1 \warp_pool_wr_data_out_reg[24]  ( .D(n773), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[24]), .QN(n92) );
  DFFR_X1 \warp_pool_wr_data_out_reg[23]  ( .D(n774), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[23]), .QN(n93) );
  DFFR_X1 \warp_pool_wr_data_out_reg[22]  ( .D(n775), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[22]), .QN(n94) );
  DFFR_X1 \warp_pool_wr_data_out_reg[21]  ( .D(n776), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[21]), .QN(n95) );
  DFFR_X1 \warp_pool_wr_data_out_reg[20]  ( .D(n777), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[20]), .QN(n96) );
  DFFR_X1 \warp_pool_wr_data_out_reg[19]  ( .D(n778), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[19]), .QN(n97) );
  DFFR_X1 \warp_pool_wr_data_out_reg[18]  ( .D(n779), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[18]), .QN(n98) );
  DFFR_X1 \warp_pool_wr_data_out_reg[17]  ( .D(n780), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[17]), .QN(n99) );
  DFFR_X1 \warp_pool_wr_data_out_reg[16]  ( .D(n781), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[16]), .QN(n100) );
  DFFR_X1 \warp_pool_wr_data_out_reg[15]  ( .D(n782), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[15]), .QN(n101) );
  DFFR_X1 \warp_pool_wr_data_out_reg[14]  ( .D(n783), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[14]), .QN(n102) );
  DFFR_X1 \warp_pool_wr_data_out_reg[13]  ( .D(n784), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[13]), .QN(n103) );
  DFFR_X1 \warp_pool_wr_data_out_reg[12]  ( .D(n785), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[12]), .QN(n104) );
  DFFR_X1 \warp_pool_wr_data_out_reg[11]  ( .D(n786), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[11]), .QN(n105) );
  DFFR_X1 \warp_pool_wr_data_out_reg[10]  ( .D(n787), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[10]), .QN(n106) );
  DFFR_X1 \warp_pool_wr_data_out_reg[9]  ( .D(n788), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[9]), .QN(n107) );
  DFFR_X1 \warp_pool_wr_data_out_reg[8]  ( .D(n789), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[8]), .QN(n108) );
  DFFR_X1 \warp_pool_wr_data_out_reg[7]  ( .D(n790), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[7]), .QN(n109) );
  DFFR_X1 \warp_pool_wr_data_out_reg[6]  ( .D(n791), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[6]), .QN(n110) );
  DFFR_X1 \warp_pool_wr_data_out_reg[5]  ( .D(n792), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[5]), .QN(n111) );
  DFFR_X1 \warp_pool_wr_data_out_reg[4]  ( .D(n793), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[4]), .QN(n112) );
  DFFR_X1 \warp_pool_wr_data_out_reg[3]  ( .D(n794), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[3]), .QN(n113) );
  DFFR_X1 \warp_pool_wr_data_out_reg[2]  ( .D(n795), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[2]), .QN(n114) );
  DFFR_X1 \warp_pool_wr_data_out_reg[1]  ( .D(n796), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[1]), .QN(n115) );
  DFFR_X1 \warp_num_i_reg[0]  ( .D(n802), .CK(clk_in), .RN(n125), .Q(
        warp_num_i[0]) );
  DFFR_X1 \warp_num_i_reg[1]  ( .D(n803), .CK(clk_in), .RN(n125), .Q(
        warp_num_i[1]) );
  DFFR_X1 \warp_num_i_reg[2]  ( .D(n804), .CK(clk_in), .RN(n125), .Q(
        warp_num_i[2]) );
  DFFR_X1 \warp_num_i_reg[3]  ( .D(n805), .CK(clk_in), .RN(n125), .Q(
        warp_num_i[3]) );
  DFFR_X1 \warp_num_i_reg[4]  ( .D(n806), .CK(clk_in), .RN(n125), .Q(
        warp_num_i[4]) );
  DFFR_X1 warp_id_calc_en_i_reg ( .D(n798), .CK(clk_in), .RN(n125), .Q(
        warp_id_calc_en_i), .QN(n156) );
  DFFR_X1 \block_num_i_reg[1]  ( .D(n799), .CK(clk_in), .RN(n125), .Q(
        block_num_i[1]), .QN(n154) );
  DFFR_X1 \warp_pool_wr_data_out_reg[107]  ( .D(n731), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[107]), .QN(n42) );
  DFFR_X1 \block_num_i_reg[2]  ( .D(n800), .CK(clk_in), .RN(n125), .Q(
        block_num_i[2]), .QN(n153) );
  DFFR_X1 \warp_pool_wr_data_out_reg[108]  ( .D(n730), .CK(clk_in), .RN(n126), 
        .Q(warp_pool_wr_data_out[108]), .QN(n41) );
  DFFR_X1 \block_num_i_reg[3]  ( .D(n801), .CK(clk_in), .RN(n126), .Q(
        block_num_i[3]), .QN(n152) );
  DFFR_X1 \warp_pool_wr_data_out_reg[109]  ( .D(n729), .CK(clk_in), .RN(n126), 
        .Q(warp_pool_wr_data_out[109]), .QN(n40) );
  DFFR_X1 \block_num_i_reg[0]  ( .D(n807), .CK(clk_in), .RN(n126), .Q(
        block_num_i[0]), .QN(n155) );
  DFFR_X1 \warp_state_addr_out_reg[0]  ( .D(n182), .CK(clk_in), .RN(n126), .Q(
        warp_state_addr_out[0]) );
  DFFR_X1 \warp_pool_addr_out_reg[0]  ( .D(n181), .CK(clk_in), .RN(n126), .Q(
        warp_pool_addr_out[0]) );
  DFFR_X1 \warp_state_addr_out_reg[1]  ( .D(n177), .CK(clk_in), .RN(n126), .Q(
        warp_state_addr_out[1]) );
  DFFR_X1 \warp_pool_addr_out_reg[1]  ( .D(n176), .CK(clk_in), .RN(n126), .Q(
        warp_pool_addr_out[1]) );
  DFFR_X1 \warp_state_addr_out_reg[2]  ( .D(n173), .CK(clk_in), .RN(n126), .Q(
        warp_state_addr_out[2]) );
  DFFR_X1 \warp_pool_addr_out_reg[2]  ( .D(n172), .CK(clk_in), .RN(n126), .Q(
        warp_pool_addr_out[2]) );
  DFFR_X1 \warp_state_addr_out_reg[3]  ( .D(n169), .CK(clk_in), .RN(n126), .Q(
        warp_state_addr_out[3]) );
  DFFR_X1 \warp_pool_addr_out_reg[3]  ( .D(n168), .CK(clk_in), .RN(n126), .Q(
        warp_pool_addr_out[3]) );
  DFFR_X1 \warp_state_addr_out_reg[4]  ( .D(n165), .CK(clk_in), .RN(n126), .Q(
        warp_state_addr_out[4]) );
  DFFR_X1 \warp_pool_addr_out_reg[4]  ( .D(n164), .CK(clk_in), .RN(n126), .Q(
        warp_pool_addr_out[4]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[97]  ( .D(n178), .CK(clk_in), .RN(n126), 
        .Q(warp_pool_wr_data_out[97]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[98]  ( .D(n161), .CK(clk_in), .RN(n126), 
        .Q(warp_pool_wr_data_out[98]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[99]  ( .D(n160), .CK(clk_in), .RN(n126), 
        .Q(warp_pool_wr_data_out[99]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[100]  ( .D(n159), .CK(clk_in), .RN(n126), 
        .Q(warp_pool_wr_data_out[100]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[101]  ( .D(n158), .CK(clk_in), .RN(n126), 
        .Q(warp_pool_wr_data_out[101]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[102]  ( .D(n157), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[102]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[103]  ( .D(n146), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[103]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[104]  ( .D(n144), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[104]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[105]  ( .D(n140), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[105]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[106]  ( .D(n732), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[106]), .QN(n43) );
  DFFR_X1 warp_gen_done_reg ( .D(n797), .CK(clk_in), .RN(n127), .Q(
        warp_gen_done) );
  DFFR_X1 \num_warps_out_reg[1]  ( .D(n174), .CK(clk_in), .RN(n127), .Q(
        num_warps_out[1]) );
  DFFR_X1 \num_warps_out_reg[2]  ( .D(n170), .CK(clk_in), .RN(n127), .Q(
        num_warps_out[2]) );
  DFFR_X1 \num_warps_out_reg[3]  ( .D(n166), .CK(clk_in), .RN(n127), .Q(
        num_warps_out[3]) );
  DFFR_X1 \num_warps_out_reg[4]  ( .D(n162), .CK(clk_in), .RN(n127), .Q(
        num_warps_out[4]) );
  DFFR_X1 \num_warps_out_reg[0]  ( .D(n179), .CK(clk_in), .RN(n127), .Q(
        num_warps_out[0]) );
  DFF_X1 \shmem_addr_i_reg[13]  ( .D(n183), .CK(clk_in), .Q(shmem_addr_i[13])
         );
  DFFR_X1 \warp_pool_wr_data_out_reg[123]  ( .D(n858), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[123]) );
  DFF_X1 \shmem_addr_i_reg[12]  ( .D(n184), .CK(clk_in), .Q(shmem_addr_i[12])
         );
  DFFR_X1 \warp_pool_wr_data_out_reg[122]  ( .D(n859), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[122]) );
  DFF_X1 \shmem_addr_i_reg[11]  ( .D(n185), .CK(clk_in), .Q(shmem_addr_i[11])
         );
  DFFR_X1 \warp_pool_wr_data_out_reg[121]  ( .D(n860), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[121]) );
  DFF_X1 \shmem_addr_i_reg[10]  ( .D(n186), .CK(clk_in), .Q(shmem_addr_i[10])
         );
  DFFR_X1 \warp_pool_wr_data_out_reg[120]  ( .D(n861), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[120]) );
  DFF_X1 \shmem_addr_i_reg[9]  ( .D(n187), .CK(clk_in), .Q(shmem_addr_i[9]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[119]  ( .D(n862), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[119]) );
  DFF_X1 \shmem_addr_i_reg[8]  ( .D(n188), .CK(clk_in), .Q(shmem_addr_i[8]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[118]  ( .D(n863), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[118]) );
  DFF_X1 \shmem_addr_i_reg[7]  ( .D(n189), .CK(clk_in), .Q(shmem_addr_i[7]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[117]  ( .D(n864), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[117]) );
  DFF_X1 \shmem_addr_i_reg[6]  ( .D(n190), .CK(clk_in), .Q(shmem_addr_i[6]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[116]  ( .D(n865), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[116]) );
  DFF_X1 \shmem_addr_i_reg[5]  ( .D(n191), .CK(clk_in), .Q(shmem_addr_i[5]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[115]  ( .D(n866), .CK(clk_in), .RN(n127), 
        .Q(warp_pool_wr_data_out[115]) );
  DFF_X1 \shmem_addr_i_reg[4]  ( .D(n192), .CK(clk_in), .Q(shmem_addr_i[4]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[114]  ( .D(n867), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[114]) );
  DFF_X1 \shmem_addr_i_reg[3]  ( .D(n193), .CK(clk_in), .Q(shmem_addr_i[3]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[113]  ( .D(n868), .CK(clk_in), .RN(n123), 
        .Q(warp_pool_wr_data_out[113]) );
  DFF_X1 \shmem_addr_i_reg[2]  ( .D(n194), .CK(clk_in), .Q(shmem_addr_i[2]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[112]  ( .D(n869), .CK(clk_in), .RN(n124), 
        .Q(warp_pool_wr_data_out[112]) );
  DFF_X1 \shmem_addr_i_reg[1]  ( .D(n195), .CK(clk_in), .Q(shmem_addr_i[1]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[111]  ( .D(n870), .CK(clk_in), .RN(n125), 
        .Q(warp_pool_wr_data_out[111]) );
  DFF_X1 \shmem_addr_i_reg[0]  ( .D(n196), .CK(clk_in), .Q(shmem_addr_i[0]) );
  DFFR_X1 \warp_pool_wr_data_out_reg[110]  ( .D(n871), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[110]) );
  DFF_X1 \warp_id_addr_reg[4]  ( .D(n728), .CK(clk_in), .Q(warp_id_addr[4]), 
        .QN(n267) );
  DFF_X1 \warp_id_addr_reg[3]  ( .D(n727), .CK(clk_in), .Q(warp_id_addr[3]), 
        .QN(n268) );
  DFF_X1 \warp_id_addr_reg[2]  ( .D(n726), .CK(clk_in), .Q(warp_id_addr[2]), 
        .QN(n269) );
  DFF_X1 \warp_id_addr_reg[1]  ( .D(n725), .CK(clk_in), .Q(warp_id_addr[1]), 
        .QN(n270) );
  DFF_X1 \warp_id_addr_reg[0]  ( .D(n724), .CK(clk_in), .Q(warp_id_addr[0]), 
        .QN(n271) );
  DFF_X1 \fence_regs_cta_id_out_reg[25><3]  ( .D(n620), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[25><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[25><2]  ( .D(n621), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[25><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[25><1]  ( .D(n622), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[25><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[25><0]  ( .D(n623), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[25><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[25]  ( .D(n538), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[25]), .QN(n241) );
  DFF_X1 \fence_regs_cta_id_ld_reg[25]  ( .D(n570), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[25]), .QN(n209) );
  DFF_X1 \fence_regs_cta_id_out_reg[17><3]  ( .D(n652), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[17><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[17><2]  ( .D(n653), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[17><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[17><1]  ( .D(n654), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[17><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[17><0]  ( .D(n655), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[17><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[17]  ( .D(n546), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[17]), .QN(n249) );
  DFF_X1 \fence_regs_cta_id_ld_reg[17]  ( .D(n578), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[17]), .QN(n217) );
  DFF_X1 \fence_regs_cta_id_out_reg[9><3]  ( .D(n684), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[9><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[9><2]  ( .D(n685), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[9><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[9><1]  ( .D(n686), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[9><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[9><0]  ( .D(n687), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[9><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[9]  ( .D(n554), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[9]), .QN(n257) );
  DFF_X1 \fence_regs_cta_id_ld_reg[9]  ( .D(n586), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[9]), .QN(n225) );
  DFF_X1 \fence_regs_cta_id_out_reg[1><3]  ( .D(n716), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[1><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[1><2]  ( .D(n717), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[1><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[1><1]  ( .D(n718), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[1><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[1><0]  ( .D(n719), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[1><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[1]  ( .D(n562), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[1]), .QN(n265) );
  DFF_X1 \fence_regs_cta_id_ld_reg[1]  ( .D(n594), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[1]), .QN(n233) );
  DFF_X1 \fence_regs_cta_id_out_reg[27><3]  ( .D(n612), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[27><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[27><2]  ( .D(n613), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[27><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[27><1]  ( .D(n614), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[27><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[27><0]  ( .D(n615), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[27><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[27]  ( .D(n536), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[27]), .QN(n239) );
  DFF_X1 \fence_regs_cta_id_ld_reg[27]  ( .D(n568), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[27]), .QN(n207) );
  DFF_X1 \fence_regs_cta_id_out_reg[19><3]  ( .D(n644), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[19><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[19><2]  ( .D(n645), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[19><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[19><1]  ( .D(n646), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[19><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[19><0]  ( .D(n647), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[19><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[19]  ( .D(n544), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[19]), .QN(n247) );
  DFF_X1 \fence_regs_cta_id_ld_reg[19]  ( .D(n576), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[19]), .QN(n215) );
  DFF_X1 \fence_regs_cta_id_out_reg[11><3]  ( .D(n676), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[11><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[11><2]  ( .D(n677), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[11><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[11><1]  ( .D(n678), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[11><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[11><0]  ( .D(n679), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[11><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[11]  ( .D(n552), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[11]), .QN(n255) );
  DFF_X1 \fence_regs_cta_id_ld_reg[11]  ( .D(n584), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[11]), .QN(n223) );
  DFF_X1 \fence_regs_cta_id_out_reg[3><3]  ( .D(n708), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[3><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[3><2]  ( .D(n709), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[3><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[3><1]  ( .D(n710), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[3><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[3><0]  ( .D(n711), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[3><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[3]  ( .D(n560), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[3]), .QN(n263) );
  DFF_X1 \fence_regs_cta_id_ld_reg[3]  ( .D(n592), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[3]), .QN(n231) );
  DFF_X1 \fence_regs_cta_id_out_reg[29><3]  ( .D(n604), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[29><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[29><2]  ( .D(n605), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[29><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[29><1]  ( .D(n606), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[29><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[29><0]  ( .D(n607), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[29><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[29]  ( .D(n534), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[29]), .QN(n237) );
  DFF_X1 \fence_regs_cta_id_ld_reg[29]  ( .D(n566), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[29]), .QN(n205) );
  DFF_X1 \fence_regs_cta_id_out_reg[21><3]  ( .D(n636), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[21><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[21><2]  ( .D(n637), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[21><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[21><1]  ( .D(n638), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[21><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[21><0]  ( .D(n639), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[21><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[21]  ( .D(n542), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[21]), .QN(n245) );
  DFF_X1 \fence_regs_cta_id_ld_reg[21]  ( .D(n574), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[21]), .QN(n213) );
  DFF_X1 \fence_regs_cta_id_out_reg[13><3]  ( .D(n668), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[13><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[13><2]  ( .D(n669), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[13><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[13><1]  ( .D(n670), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[13><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[13><0]  ( .D(n671), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[13><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[13]  ( .D(n550), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[13]), .QN(n253) );
  DFF_X1 \fence_regs_cta_id_ld_reg[13]  ( .D(n582), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[13]), .QN(n221) );
  DFF_X1 \fence_regs_cta_id_out_reg[5><3]  ( .D(n700), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[5><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[5><2]  ( .D(n701), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[5><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[5><1]  ( .D(n702), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[5><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[5><0]  ( .D(n703), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[5><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[5]  ( .D(n558), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[5]), .QN(n261) );
  DFF_X1 \fence_regs_cta_id_ld_reg[5]  ( .D(n590), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[5]), .QN(n229) );
  DFF_X1 \fence_regs_cta_id_out_reg[31><3]  ( .D(n596), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[31><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[31><2]  ( .D(n597), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[31><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[31><1]  ( .D(n598), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[31><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[31><0]  ( .D(n599), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[31><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[31]  ( .D(n532), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[31]), .QN(n235) );
  DFF_X1 \fence_regs_cta_id_ld_reg[31]  ( .D(n564), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[31]), .QN(n203) );
  DFF_X1 \fence_regs_cta_id_out_reg[23><3]  ( .D(n628), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[23><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[23><2]  ( .D(n629), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[23><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[23><1]  ( .D(n630), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[23><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[23><0]  ( .D(n631), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[23><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[23]  ( .D(n540), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[23]), .QN(n243) );
  DFF_X1 \fence_regs_cta_id_ld_reg[23]  ( .D(n572), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[23]), .QN(n211) );
  DFF_X1 \fence_regs_cta_id_out_reg[15><3]  ( .D(n660), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[15><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[15><2]  ( .D(n661), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[15><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[15><1]  ( .D(n662), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[15><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[15><0]  ( .D(n663), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[15><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[15]  ( .D(n548), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[15]), .QN(n251) );
  DFF_X1 \fence_regs_cta_id_ld_reg[15]  ( .D(n580), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[15]), .QN(n219) );
  DFF_X1 \fence_regs_cta_id_out_reg[7><3]  ( .D(n692), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[7><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[7><2]  ( .D(n693), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[7><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[7><1]  ( .D(n694), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[7><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[7><0]  ( .D(n695), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[7><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[7]  ( .D(n556), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[7]), .QN(n259) );
  DFF_X1 \fence_regs_cta_id_ld_reg[7]  ( .D(n588), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[7]), .QN(n227) );
  DFF_X1 \fence_regs_cta_id_out_reg[24><3]  ( .D(n624), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[24><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[24><2]  ( .D(n625), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[24><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[24><1]  ( .D(n626), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[24><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[24><0]  ( .D(n627), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[24><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[24]  ( .D(n539), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[24]), .QN(n242) );
  DFF_X1 \fence_regs_cta_id_ld_reg[24]  ( .D(n571), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[24]), .QN(n210) );
  DFF_X1 \fence_regs_cta_id_out_reg[16><3]  ( .D(n656), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[16><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[16><2]  ( .D(n657), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[16><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[16><1]  ( .D(n658), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[16><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[16><0]  ( .D(n659), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[16><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[16]  ( .D(n547), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[16]), .QN(n250) );
  DFF_X1 \fence_regs_cta_id_ld_reg[16]  ( .D(n579), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[16]), .QN(n218) );
  DFF_X1 \fence_regs_cta_id_out_reg[8><3]  ( .D(n688), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[8><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[8><2]  ( .D(n689), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[8><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[8><1]  ( .D(n690), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[8><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[8><0]  ( .D(n691), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[8><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[8]  ( .D(n555), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[8]), .QN(n258) );
  DFF_X1 \fence_regs_cta_id_ld_reg[8]  ( .D(n587), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[8]), .QN(n226) );
  DFF_X1 \fence_regs_cta_id_out_reg[0><3]  ( .D(n720), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[0><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[0><2]  ( .D(n721), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[0><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[0><1]  ( .D(n722), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[0><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[0><0]  ( .D(n723), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[0><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[0]  ( .D(n563), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[0]), .QN(n266) );
  DFF_X1 \fence_regs_cta_id_ld_reg[0]  ( .D(n595), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[0]), .QN(n234) );
  DFF_X1 \fence_regs_cta_id_out_reg[26><3]  ( .D(n616), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[26><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[26><2]  ( .D(n617), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[26><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[26><1]  ( .D(n618), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[26><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[26><0]  ( .D(n619), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[26><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[26]  ( .D(n537), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[26]), .QN(n240) );
  DFF_X1 \fence_regs_cta_id_ld_reg[26]  ( .D(n569), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[26]), .QN(n208) );
  DFF_X1 \fence_regs_cta_id_out_reg[18><3]  ( .D(n648), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[18><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[18><2]  ( .D(n649), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[18><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[18><1]  ( .D(n650), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[18><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[18><0]  ( .D(n651), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[18><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[18]  ( .D(n545), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[18]), .QN(n248) );
  DFF_X1 \fence_regs_cta_id_ld_reg[18]  ( .D(n577), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[18]), .QN(n216) );
  DFF_X1 \fence_regs_cta_id_out_reg[10><3]  ( .D(n680), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[10><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[10><2]  ( .D(n681), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[10><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[10><1]  ( .D(n682), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[10><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[10><0]  ( .D(n683), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[10><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[10]  ( .D(n553), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[10]), .QN(n256) );
  DFF_X1 \fence_regs_cta_id_ld_reg[10]  ( .D(n585), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[10]), .QN(n224) );
  DFF_X1 \fence_regs_cta_id_out_reg[2><3]  ( .D(n712), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[2><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[2><2]  ( .D(n713), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[2><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[2><1]  ( .D(n714), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[2><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[2><0]  ( .D(n715), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[2><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[2]  ( .D(n561), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[2]), .QN(n264) );
  DFF_X1 \fence_regs_cta_id_ld_reg[2]  ( .D(n593), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[2]), .QN(n232) );
  DFF_X1 \fence_regs_cta_id_out_reg[28><3]  ( .D(n608), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[28><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[28><2]  ( .D(n609), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[28><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[28><1]  ( .D(n610), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[28><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[28><0]  ( .D(n611), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[28><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[28]  ( .D(n535), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[28]), .QN(n238) );
  DFF_X1 \fence_regs_cta_id_ld_reg[28]  ( .D(n567), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[28]), .QN(n206) );
  DFF_X1 \fence_regs_cta_id_out_reg[20><3]  ( .D(n640), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[20><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[20><2]  ( .D(n641), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[20><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[20><1]  ( .D(n642), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[20><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[20><0]  ( .D(n643), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[20><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[20]  ( .D(n543), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[20]), .QN(n246) );
  DFF_X1 \fence_regs_cta_id_ld_reg[20]  ( .D(n575), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[20]), .QN(n214) );
  DFF_X1 \fence_regs_cta_id_out_reg[12><3]  ( .D(n672), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[12><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[12><2]  ( .D(n673), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[12><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[12><1]  ( .D(n674), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[12><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[12><0]  ( .D(n675), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[12><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[12]  ( .D(n551), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[12]), .QN(n254) );
  DFF_X1 \fence_regs_cta_id_ld_reg[12]  ( .D(n583), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[12]), .QN(n222) );
  DFF_X1 \fence_regs_cta_id_out_reg[4><3]  ( .D(n704), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[4><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[4><2]  ( .D(n705), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[4><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[4><1]  ( .D(n706), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[4><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[4><0]  ( .D(n707), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[4><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[4]  ( .D(n559), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[4]), .QN(n262) );
  DFF_X1 \fence_regs_cta_id_ld_reg[4]  ( .D(n591), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[4]), .QN(n230) );
  DFF_X1 \fence_regs_cta_id_out_reg[30><3]  ( .D(n600), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[30><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[30><2]  ( .D(n601), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[30><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[30><1]  ( .D(n602), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[30><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[30><0]  ( .D(n603), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[30><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[30]  ( .D(n533), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[30]), .QN(n236) );
  DFF_X1 \fence_regs_cta_id_ld_reg[30]  ( .D(n565), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[30]), .QN(n204) );
  DFF_X1 \fence_regs_cta_id_out_reg[22><3]  ( .D(n632), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[22><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[22><2]  ( .D(n633), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[22><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[22><1]  ( .D(n634), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[22><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[22><0]  ( .D(n635), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[22><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[22]  ( .D(n541), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[22]), .QN(n244) );
  DFF_X1 \fence_regs_cta_id_ld_reg[22]  ( .D(n573), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[22]), .QN(n212) );
  DFF_X1 \fence_regs_cta_id_out_reg[14><3]  ( .D(n664), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[14><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[14><2]  ( .D(n665), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[14><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[14><1]  ( .D(n666), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[14><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[14><0]  ( .D(n667), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[14><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[14]  ( .D(n549), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[14]), .QN(n252) );
  DFF_X1 \fence_regs_cta_id_ld_reg[14]  ( .D(n581), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[14]), .QN(n220) );
  DFF_X1 \fence_regs_cta_id_out_reg[6><3]  ( .D(n696), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[6><3] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[6><2]  ( .D(n697), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[6><2] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[6><1]  ( .D(n698), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[6><1] ) );
  DFF_X1 \fence_regs_cta_id_out_reg[6><0]  ( .D(n699), .CK(clk_in), .Q(
        \fence_regs_cta_id_out[6><0] ) );
  DFF_X1 \fence_regs_fence_en_ld_reg[6]  ( .D(n557), .CK(clk_in), .Q(
        fence_regs_fence_en_ld[6]), .QN(n260) );
  DFF_X1 \fence_regs_cta_id_ld_reg[6]  ( .D(n589), .CK(clk_in), .Q(
        fence_regs_cta_id_ld[6]), .QN(n228) );
  NOR2_X2 U313 ( .A1(n439), .A2(n453), .ZN(n438) );
  NOR3_X2 U429 ( .A1(n453), .A2(n496), .A3(n873), .ZN(n495) );
  NAND2_X1 U597 ( .A1(\fence_regs_cta_id_out[31><3] ), .A2(n856), .ZN(n281) );
  NAND2_X1 U598 ( .A1(\fence_regs_cta_id_out[31><2] ), .A2(n856), .ZN(n283) );
  NAND2_X1 U599 ( .A1(\fence_regs_cta_id_out[31><1] ), .A2(n856), .ZN(n285) );
  NAND2_X1 U600 ( .A1(\fence_regs_cta_id_out[31><0] ), .A2(n856), .ZN(n287) );
  NAND2_X1 U601 ( .A1(\fence_regs_cta_id_out[30><3] ), .A2(n855), .ZN(n288) );
  NAND2_X1 U602 ( .A1(\fence_regs_cta_id_out[30><2] ), .A2(n855), .ZN(n289) );
  NAND2_X1 U603 ( .A1(\fence_regs_cta_id_out[30><1] ), .A2(n855), .ZN(n290) );
  NAND2_X1 U604 ( .A1(\fence_regs_cta_id_out[30><0] ), .A2(n855), .ZN(n291) );
  NAND2_X1 U605 ( .A1(\fence_regs_cta_id_out[29><3] ), .A2(n854), .ZN(n292) );
  NAND2_X1 U606 ( .A1(\fence_regs_cta_id_out[29><2] ), .A2(n854), .ZN(n293) );
  NAND2_X1 U607 ( .A1(\fence_regs_cta_id_out[29><1] ), .A2(n854), .ZN(n294) );
  NAND2_X1 U608 ( .A1(\fence_regs_cta_id_out[29><0] ), .A2(n854), .ZN(n295) );
  NAND2_X1 U609 ( .A1(\fence_regs_cta_id_out[28><3] ), .A2(n853), .ZN(n296) );
  NAND2_X1 U610 ( .A1(\fence_regs_cta_id_out[28><2] ), .A2(n853), .ZN(n297) );
  NAND2_X1 U611 ( .A1(\fence_regs_cta_id_out[28><1] ), .A2(n853), .ZN(n298) );
  NAND2_X1 U612 ( .A1(\fence_regs_cta_id_out[28><0] ), .A2(n853), .ZN(n299) );
  NAND2_X1 U613 ( .A1(\fence_regs_cta_id_out[27><3] ), .A2(n852), .ZN(n300) );
  NAND2_X1 U614 ( .A1(\fence_regs_cta_id_out[27><2] ), .A2(n852), .ZN(n301) );
  NAND2_X1 U615 ( .A1(\fence_regs_cta_id_out[27><1] ), .A2(n852), .ZN(n302) );
  NAND2_X1 U616 ( .A1(\fence_regs_cta_id_out[27><0] ), .A2(n852), .ZN(n303) );
  NAND2_X1 U617 ( .A1(\fence_regs_cta_id_out[26><3] ), .A2(n851), .ZN(n304) );
  NAND2_X1 U618 ( .A1(\fence_regs_cta_id_out[26><2] ), .A2(n851), .ZN(n305) );
  NAND2_X1 U619 ( .A1(\fence_regs_cta_id_out[26><1] ), .A2(n851), .ZN(n306) );
  NAND2_X1 U620 ( .A1(\fence_regs_cta_id_out[26><0] ), .A2(n851), .ZN(n307) );
  NAND2_X1 U621 ( .A1(\fence_regs_cta_id_out[25><3] ), .A2(n850), .ZN(n308) );
  NAND2_X1 U622 ( .A1(\fence_regs_cta_id_out[25><2] ), .A2(n850), .ZN(n309) );
  NAND2_X1 U623 ( .A1(\fence_regs_cta_id_out[25><1] ), .A2(n850), .ZN(n310) );
  NAND2_X1 U624 ( .A1(\fence_regs_cta_id_out[25><0] ), .A2(n850), .ZN(n311) );
  NAND2_X1 U625 ( .A1(\fence_regs_cta_id_out[24><3] ), .A2(n849), .ZN(n312) );
  NAND2_X1 U626 ( .A1(\fence_regs_cta_id_out[24><2] ), .A2(n849), .ZN(n313) );
  NAND2_X1 U627 ( .A1(\fence_regs_cta_id_out[24><1] ), .A2(n849), .ZN(n314) );
  NAND2_X1 U628 ( .A1(\fence_regs_cta_id_out[24><0] ), .A2(n849), .ZN(n315) );
  NAND2_X1 U629 ( .A1(\fence_regs_cta_id_out[23><3] ), .A2(n848), .ZN(n316) );
  NAND2_X1 U630 ( .A1(\fence_regs_cta_id_out[23><2] ), .A2(n848), .ZN(n317) );
  NAND2_X1 U631 ( .A1(\fence_regs_cta_id_out[23><1] ), .A2(n848), .ZN(n318) );
  NAND2_X1 U632 ( .A1(\fence_regs_cta_id_out[23><0] ), .A2(n848), .ZN(n319) );
  NAND2_X1 U633 ( .A1(\fence_regs_cta_id_out[22><3] ), .A2(n847), .ZN(n320) );
  NAND2_X1 U634 ( .A1(\fence_regs_cta_id_out[22><2] ), .A2(n847), .ZN(n321) );
  NAND2_X1 U635 ( .A1(\fence_regs_cta_id_out[22><1] ), .A2(n847), .ZN(n322) );
  NAND2_X1 U636 ( .A1(\fence_regs_cta_id_out[22><0] ), .A2(n847), .ZN(n323) );
  NAND2_X1 U637 ( .A1(\fence_regs_cta_id_out[21><3] ), .A2(n846), .ZN(n324) );
  NAND2_X1 U638 ( .A1(\fence_regs_cta_id_out[21><2] ), .A2(n846), .ZN(n325) );
  NAND2_X1 U639 ( .A1(\fence_regs_cta_id_out[21><1] ), .A2(n846), .ZN(n326) );
  NAND2_X1 U640 ( .A1(\fence_regs_cta_id_out[21><0] ), .A2(n846), .ZN(n327) );
  NAND2_X1 U641 ( .A1(\fence_regs_cta_id_out[20><3] ), .A2(n845), .ZN(n328) );
  NAND2_X1 U642 ( .A1(\fence_regs_cta_id_out[20><2] ), .A2(n845), .ZN(n329) );
  NAND2_X1 U643 ( .A1(\fence_regs_cta_id_out[20><1] ), .A2(n845), .ZN(n330) );
  NAND2_X1 U644 ( .A1(\fence_regs_cta_id_out[20><0] ), .A2(n845), .ZN(n331) );
  NAND2_X1 U645 ( .A1(\fence_regs_cta_id_out[19><3] ), .A2(n844), .ZN(n332) );
  NAND2_X1 U646 ( .A1(\fence_regs_cta_id_out[19><2] ), .A2(n844), .ZN(n333) );
  NAND2_X1 U647 ( .A1(\fence_regs_cta_id_out[19><1] ), .A2(n844), .ZN(n334) );
  NAND2_X1 U648 ( .A1(\fence_regs_cta_id_out[19><0] ), .A2(n844), .ZN(n335) );
  NAND2_X1 U649 ( .A1(\fence_regs_cta_id_out[18><3] ), .A2(n843), .ZN(n336) );
  NAND2_X1 U650 ( .A1(\fence_regs_cta_id_out[18><2] ), .A2(n843), .ZN(n337) );
  NAND2_X1 U651 ( .A1(\fence_regs_cta_id_out[18><1] ), .A2(n843), .ZN(n338) );
  NAND2_X1 U652 ( .A1(\fence_regs_cta_id_out[18><0] ), .A2(n843), .ZN(n339) );
  NAND2_X1 U653 ( .A1(\fence_regs_cta_id_out[17><3] ), .A2(n842), .ZN(n340) );
  NAND2_X1 U654 ( .A1(\fence_regs_cta_id_out[17><2] ), .A2(n842), .ZN(n341) );
  NAND2_X1 U655 ( .A1(\fence_regs_cta_id_out[17><1] ), .A2(n842), .ZN(n342) );
  NAND2_X1 U656 ( .A1(\fence_regs_cta_id_out[17><0] ), .A2(n842), .ZN(n343) );
  NAND2_X1 U657 ( .A1(\fence_regs_cta_id_out[16><3] ), .A2(n841), .ZN(n344) );
  NAND2_X1 U658 ( .A1(\fence_regs_cta_id_out[16><2] ), .A2(n841), .ZN(n345) );
  NAND2_X1 U659 ( .A1(\fence_regs_cta_id_out[16><1] ), .A2(n841), .ZN(n346) );
  NAND2_X1 U660 ( .A1(\fence_regs_cta_id_out[16><0] ), .A2(n841), .ZN(n347) );
  NAND2_X1 U661 ( .A1(\fence_regs_cta_id_out[15><3] ), .A2(n840), .ZN(n348) );
  NAND2_X1 U662 ( .A1(\fence_regs_cta_id_out[15><2] ), .A2(n840), .ZN(n349) );
  NAND2_X1 U663 ( .A1(\fence_regs_cta_id_out[15><1] ), .A2(n840), .ZN(n350) );
  NAND2_X1 U664 ( .A1(\fence_regs_cta_id_out[15><0] ), .A2(n840), .ZN(n351) );
  NAND2_X1 U665 ( .A1(\fence_regs_cta_id_out[14><3] ), .A2(n839), .ZN(n352) );
  NAND2_X1 U666 ( .A1(\fence_regs_cta_id_out[14><2] ), .A2(n839), .ZN(n353) );
  NAND2_X1 U667 ( .A1(\fence_regs_cta_id_out[14><1] ), .A2(n839), .ZN(n354) );
  NAND2_X1 U668 ( .A1(\fence_regs_cta_id_out[14><0] ), .A2(n839), .ZN(n355) );
  NAND2_X1 U669 ( .A1(\fence_regs_cta_id_out[13><3] ), .A2(n838), .ZN(n356) );
  NAND2_X1 U670 ( .A1(\fence_regs_cta_id_out[13><2] ), .A2(n838), .ZN(n357) );
  NAND2_X1 U671 ( .A1(\fence_regs_cta_id_out[13><1] ), .A2(n838), .ZN(n358) );
  NAND2_X1 U672 ( .A1(\fence_regs_cta_id_out[13><0] ), .A2(n838), .ZN(n359) );
  NAND2_X1 U673 ( .A1(\fence_regs_cta_id_out[12><3] ), .A2(n837), .ZN(n360) );
  NAND2_X1 U674 ( .A1(\fence_regs_cta_id_out[12><2] ), .A2(n837), .ZN(n361) );
  NAND2_X1 U675 ( .A1(\fence_regs_cta_id_out[12><1] ), .A2(n837), .ZN(n362) );
  NAND2_X1 U676 ( .A1(\fence_regs_cta_id_out[12><0] ), .A2(n837), .ZN(n363) );
  NAND2_X1 U677 ( .A1(\fence_regs_cta_id_out[11><3] ), .A2(n836), .ZN(n364) );
  NAND2_X1 U678 ( .A1(\fence_regs_cta_id_out[11><2] ), .A2(n836), .ZN(n365) );
  NAND2_X1 U679 ( .A1(\fence_regs_cta_id_out[11><1] ), .A2(n836), .ZN(n366) );
  NAND2_X1 U680 ( .A1(\fence_regs_cta_id_out[11><0] ), .A2(n836), .ZN(n367) );
  NAND2_X1 U681 ( .A1(\fence_regs_cta_id_out[10><3] ), .A2(n835), .ZN(n368) );
  NAND2_X1 U682 ( .A1(\fence_regs_cta_id_out[10><2] ), .A2(n835), .ZN(n369) );
  NAND2_X1 U683 ( .A1(\fence_regs_cta_id_out[10><1] ), .A2(n835), .ZN(n370) );
  NAND2_X1 U684 ( .A1(\fence_regs_cta_id_out[10><0] ), .A2(n835), .ZN(n371) );
  NAND2_X1 U685 ( .A1(\fence_regs_cta_id_out[9><3] ), .A2(n834), .ZN(n372) );
  NAND2_X1 U686 ( .A1(\fence_regs_cta_id_out[9><2] ), .A2(n834), .ZN(n373) );
  NAND2_X1 U687 ( .A1(\fence_regs_cta_id_out[9><1] ), .A2(n834), .ZN(n374) );
  NAND2_X1 U688 ( .A1(\fence_regs_cta_id_out[9><0] ), .A2(n834), .ZN(n375) );
  NAND2_X1 U689 ( .A1(\fence_regs_cta_id_out[8><3] ), .A2(n833), .ZN(n376) );
  NAND2_X1 U690 ( .A1(\fence_regs_cta_id_out[8><2] ), .A2(n833), .ZN(n377) );
  NAND2_X1 U691 ( .A1(\fence_regs_cta_id_out[8><1] ), .A2(n833), .ZN(n378) );
  NAND2_X1 U692 ( .A1(\fence_regs_cta_id_out[8><0] ), .A2(n833), .ZN(n379) );
  NAND2_X1 U693 ( .A1(\fence_regs_cta_id_out[7><3] ), .A2(n832), .ZN(n380) );
  NAND2_X1 U694 ( .A1(\fence_regs_cta_id_out[7><2] ), .A2(n832), .ZN(n381) );
  NAND2_X1 U695 ( .A1(\fence_regs_cta_id_out[7><1] ), .A2(n832), .ZN(n382) );
  NAND2_X1 U696 ( .A1(\fence_regs_cta_id_out[7><0] ), .A2(n832), .ZN(n383) );
  NAND2_X1 U697 ( .A1(\fence_regs_cta_id_out[6><3] ), .A2(n831), .ZN(n384) );
  NAND2_X1 U698 ( .A1(\fence_regs_cta_id_out[6><2] ), .A2(n831), .ZN(n385) );
  NAND2_X1 U699 ( .A1(\fence_regs_cta_id_out[6><1] ), .A2(n831), .ZN(n386) );
  NAND2_X1 U700 ( .A1(\fence_regs_cta_id_out[6><0] ), .A2(n831), .ZN(n387) );
  NAND2_X1 U701 ( .A1(\fence_regs_cta_id_out[5><3] ), .A2(n830), .ZN(n388) );
  NAND2_X1 U702 ( .A1(\fence_regs_cta_id_out[5><2] ), .A2(n830), .ZN(n389) );
  NAND2_X1 U703 ( .A1(\fence_regs_cta_id_out[5><1] ), .A2(n830), .ZN(n390) );
  NAND2_X1 U704 ( .A1(\fence_regs_cta_id_out[5><0] ), .A2(n830), .ZN(n391) );
  NAND2_X1 U705 ( .A1(\fence_regs_cta_id_out[4><3] ), .A2(n829), .ZN(n392) );
  NAND2_X1 U706 ( .A1(\fence_regs_cta_id_out[4><2] ), .A2(n829), .ZN(n393) );
  NAND2_X1 U707 ( .A1(\fence_regs_cta_id_out[4><1] ), .A2(n829), .ZN(n394) );
  NAND2_X1 U708 ( .A1(\fence_regs_cta_id_out[4><0] ), .A2(n829), .ZN(n395) );
  NAND2_X1 U709 ( .A1(\fence_regs_cta_id_out[3><3] ), .A2(n828), .ZN(n396) );
  NAND2_X1 U710 ( .A1(\fence_regs_cta_id_out[3><2] ), .A2(n828), .ZN(n397) );
  NAND2_X1 U711 ( .A1(\fence_regs_cta_id_out[3><1] ), .A2(n828), .ZN(n398) );
  NAND2_X1 U712 ( .A1(\fence_regs_cta_id_out[3><0] ), .A2(n828), .ZN(n399) );
  NAND2_X1 U713 ( .A1(\fence_regs_cta_id_out[2><3] ), .A2(n827), .ZN(n400) );
  NAND2_X1 U714 ( .A1(\fence_regs_cta_id_out[2><2] ), .A2(n827), .ZN(n401) );
  NAND2_X1 U715 ( .A1(\fence_regs_cta_id_out[2><1] ), .A2(n827), .ZN(n402) );
  NAND2_X1 U716 ( .A1(\fence_regs_cta_id_out[2><0] ), .A2(n827), .ZN(n403) );
  NAND2_X1 U717 ( .A1(\fence_regs_cta_id_out[1><3] ), .A2(n826), .ZN(n404) );
  NAND2_X1 U718 ( .A1(\fence_regs_cta_id_out[1><2] ), .A2(n826), .ZN(n405) );
  NAND2_X1 U719 ( .A1(\fence_regs_cta_id_out[1><1] ), .A2(n826), .ZN(n406) );
  NAND2_X1 U720 ( .A1(\fence_regs_cta_id_out[1><0] ), .A2(n826), .ZN(n407) );
  NAND2_X1 U721 ( .A1(\fence_regs_cta_id_out[0><3] ), .A2(n825), .ZN(n408) );
  NAND2_X1 U722 ( .A1(block_num_i[3]), .A2(n34), .ZN(n280) );
  NAND2_X1 U723 ( .A1(\fence_regs_cta_id_out[0><2] ), .A2(n825), .ZN(n409) );
  NAND2_X1 U724 ( .A1(block_num_i[2]), .A2(n34), .ZN(n282) );
  NAND2_X1 U725 ( .A1(\fence_regs_cta_id_out[0><1] ), .A2(n825), .ZN(n410) );
  NAND2_X1 U726 ( .A1(block_num_i[1]), .A2(n35), .ZN(n284) );
  NAND2_X1 U727 ( .A1(\fence_regs_cta_id_out[0><0] ), .A2(n825), .ZN(n411) );
  NAND2_X1 U728 ( .A1(block_num_i[0]), .A2(n35), .ZN(n286) );
  NAND2_X1 U731 ( .A1(n455), .A2(n460), .ZN(n797) );
  NAND2_X1 U732 ( .A1(warp_gen_done), .A2(n461), .ZN(n460) );
  NAND2_X1 U733 ( .A1(warp_num_i[0]), .A2(n475), .ZN(n474) );
  NAND2_X1 U734 ( .A1(warp_num_i[1]), .A2(n475), .ZN(n476) );
  NAND2_X1 U735 ( .A1(warp_num_i[2]), .A2(n475), .ZN(n477) );
  NAND2_X1 U736 ( .A1(warp_num_i[3]), .A2(n475), .ZN(n478) );
  NAND2_X1 U737 ( .A1(warp_num_i[4]), .A2(n475), .ZN(n479) );
  NAND2_X1 U738 ( .A1(n872), .A2(n274), .ZN(n473) );
  NAND2_X1 U739 ( .A1(block_num_cnt[1]), .A2(n142), .ZN(n485) );
  NAND3_X1 U740 ( .A1(n275), .A2(n145), .A3(n872), .ZN(n487) );
  NAND3_X1 U741 ( .A1(n872), .A2(n275), .A3(block_num_cnt[0]), .ZN(n483) );
  NAND2_X1 U742 ( .A1(n489), .A2(n22), .ZN(n812) );
  NAND2_X1 U743 ( .A1(warp_state_wr_en_out), .A2(n490), .ZN(n489) );
  NAND2_X1 U744 ( .A1(n491), .A2(n22), .ZN(n813) );
  NAND2_X1 U745 ( .A1(warp_pool_wr_en_out), .A2(n490), .ZN(n491) );
  NAND3_X1 U746 ( .A1(n202), .A2(n201), .A3(warp_generator_state_machine[2]), 
        .ZN(n455) );
  NAND3_X1 U747 ( .A1(warp_id_addr[3]), .A2(n528), .A3(warp_id_addr[4]), .ZN(
        n518) );
  NAND3_X1 U748 ( .A1(n528), .A2(n268), .A3(warp_id_addr[4]), .ZN(n529) );
  NAND3_X1 U749 ( .A1(n528), .A2(n267), .A3(warp_id_addr[3]), .ZN(n530) );
  NAND3_X1 U750 ( .A1(warp_id_addr[1]), .A2(warp_id_addr[0]), .A3(
        warp_id_addr[2]), .ZN(n519) );
  NAND3_X1 U751 ( .A1(warp_id_addr[1]), .A2(n271), .A3(warp_id_addr[2]), .ZN(
        n521) );
  NAND3_X1 U752 ( .A1(warp_id_addr[0]), .A2(n270), .A3(warp_id_addr[2]), .ZN(
        n522) );
  NAND3_X1 U753 ( .A1(n271), .A2(n270), .A3(warp_id_addr[2]), .ZN(n523) );
  NAND3_X1 U754 ( .A1(warp_id_addr[0]), .A2(n269), .A3(warp_id_addr[1]), .ZN(
        n524) );
  NAND3_X1 U755 ( .A1(n271), .A2(n269), .A3(warp_id_addr[1]), .ZN(n525) );
  NAND3_X1 U756 ( .A1(n270), .A2(n269), .A3(warp_id_addr[0]), .ZN(n526) );
  NAND3_X1 U757 ( .A1(n201), .A2(n200), .A3(warp_generator_state_machine[0]), 
        .ZN(n453) );
  NAND3_X1 U758 ( .A1(n268), .A2(n267), .A3(n528), .ZN(n531) );
  NAND3_X1 U759 ( .A1(n270), .A2(n269), .A3(n271), .ZN(n527) );
  NAND3_X1 U762 ( .A1(n201), .A2(n200), .A3(n202), .ZN(n461) );
  warp_id_calc uWarpIdCalc ( .clk(clk_in), .reset(n119), .en(
        warp_id_calc_en_i), .block_num_in(block_num_i), .gprs_size_in(
        gprs_size_in), .warp_num_in(warp_num_i), .warps_per_block_in(
        warps_per_block_in), .gprs_base_addr_out(gprs_base_addr_o), 
        .warp_id_out(warp_id_o) );
  warp_generator_SHMEM_ADDR_SIZE14_DW01_inc_1 add_127 ( .A(warps_per_block_cnt), .SUM({N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, N93, N92}) );
  warp_generator_SHMEM_ADDR_SIZE14_DW02_mult_0 mult_124 ( .A(block_num_cnt), 
        .B(shmem_size_in[13:0]), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, N77, N76, N75, N74, N73, N72, N71, N70, N69, 
        N68, N67, N66, N65, N64}) );
  warp_generator_SHMEM_ADDR_SIZE14_DW01_add_0 add_124 ( .A(
        shmem_base_addr_in[13:0]), .B({N77, N76, N75, N74, N73, N72, N71, N70, 
        N69, N68, N67, N66, N65, N64}), .CI(1'b0), .SUM({N91, N90, N89, N88, 
        N87, N86, N85, N84, N83, N82, N81, N80, N79, N78}) );
  HA_X1 \add_155/U1_1_1  ( .A(warp_id_o[1]), .B(warp_id_o[0]), .CO(
        \add_155/carry[2] ), .S(N254) );
  HA_X1 \add_155/U1_1_2  ( .A(warp_id_o[2]), .B(\add_155/carry[2] ), .CO(
        \add_155/carry[3] ), .S(N255) );
  HA_X1 \add_155/U1_1_3  ( .A(warp_id_o[3]), .B(\add_155/carry[3] ), .CO(
        \add_155/carry[4] ), .S(N256) );
  INV_X1 U11 ( .A(n133), .ZN(n139) );
  NOR3_X1 U75 ( .A1(warp_generator_state_machine[0]), .A2(
        warp_generator_state_machine[2]), .A3(n201), .ZN(n413) );
  AND3_X1 U76 ( .A1(warp_generator_state_machine[0]), .A2(n200), .A3(
        warp_generator_state_machine[1]), .ZN(n1) );
  AND2_X1 U77 ( .A1(n461), .A2(n24), .ZN(n3) );
  INV_X1 U78 ( .A(n49), .ZN(n38) );
  INV_X1 U79 ( .A(n48), .ZN(n37) );
  INV_X1 U80 ( .A(n47), .ZN(n36) );
  NAND2_X1 U81 ( .A1(n274), .A2(n126), .ZN(n439) );
  BUF_X1 U82 ( .A(n52), .Z(n50) );
  BUF_X1 U83 ( .A(n52), .Z(n49) );
  BUF_X1 U84 ( .A(n117), .Z(n48) );
  BUF_X1 U85 ( .A(n117), .Z(n47) );
  BUF_X1 U86 ( .A(n117), .Z(n46) );
  INV_X1 U87 ( .A(n488), .ZN(n275) );
  BUF_X1 U88 ( .A(n520), .Z(n4) );
  BUF_X1 U89 ( .A(n520), .Z(n5) );
  BUF_X1 U90 ( .A(n520), .Z(n6) );
  BUF_X1 U91 ( .A(n118), .Z(n39) );
  BUF_X1 U92 ( .A(n118), .Z(n44) );
  BUF_X1 U93 ( .A(n118), .Z(n45) );
  BUF_X1 U94 ( .A(n52), .Z(n51) );
  NOR2_X2 U95 ( .A1(n857), .A2(n480), .ZN(n496) );
  INV_X1 U96 ( .A(N869), .ZN(n831) );
  INV_X1 U97 ( .A(N877), .ZN(n839) );
  INV_X1 U98 ( .A(N885), .ZN(n847) );
  INV_X1 U99 ( .A(N867), .ZN(n829) );
  INV_X1 U100 ( .A(N875), .ZN(n837) );
  INV_X1 U101 ( .A(N883), .ZN(n845) );
  INV_X1 U102 ( .A(N865), .ZN(n827) );
  INV_X1 U103 ( .A(N873), .ZN(n835) );
  INV_X1 U104 ( .A(N881), .ZN(n843) );
  INV_X1 U105 ( .A(N863), .ZN(n825) );
  INV_X1 U106 ( .A(N871), .ZN(n833) );
  INV_X1 U107 ( .A(N879), .ZN(n841) );
  INV_X1 U108 ( .A(N870), .ZN(n832) );
  INV_X1 U109 ( .A(N878), .ZN(n840) );
  INV_X1 U110 ( .A(N886), .ZN(n848) );
  INV_X1 U111 ( .A(N868), .ZN(n830) );
  INV_X1 U112 ( .A(N876), .ZN(n838) );
  INV_X1 U113 ( .A(N884), .ZN(n846) );
  INV_X1 U114 ( .A(N866), .ZN(n828) );
  INV_X1 U115 ( .A(N874), .ZN(n836) );
  INV_X1 U116 ( .A(N882), .ZN(n844) );
  INV_X1 U117 ( .A(N864), .ZN(n826) );
  INV_X1 U118 ( .A(N872), .ZN(n834) );
  INV_X1 U119 ( .A(N880), .ZN(n842) );
  INV_X1 U120 ( .A(N893), .ZN(n855) );
  INV_X1 U121 ( .A(N891), .ZN(n853) );
  INV_X1 U122 ( .A(N889), .ZN(n851) );
  INV_X1 U123 ( .A(N887), .ZN(n849) );
  INV_X1 U124 ( .A(N894), .ZN(n856) );
  INV_X1 U125 ( .A(N892), .ZN(n854) );
  INV_X1 U126 ( .A(N890), .ZN(n852) );
  INV_X1 U127 ( .A(N888), .ZN(n850) );
  INV_X1 U128 ( .A(n475), .ZN(n274) );
  AOI21_X1 U129 ( .B1(n873), .B2(n480), .A(n857), .ZN(n488) );
  NOR2_X1 U130 ( .A1(n23), .A2(n119), .ZN(n528) );
  NOR2_X1 U131 ( .A1(n872), .A2(n38), .ZN(n490) );
  BUF_X1 U132 ( .A(n3), .Z(n52) );
  BUF_X1 U133 ( .A(n3), .Z(n117) );
  INV_X1 U134 ( .A(n34), .ZN(n24) );
  INV_X1 U135 ( .A(n33), .ZN(n22) );
  INV_X1 U136 ( .A(n33), .ZN(n21) );
  INV_X1 U137 ( .A(n31), .ZN(n20) );
  INV_X1 U138 ( .A(n30), .ZN(n19) );
  INV_X1 U139 ( .A(n412), .ZN(n199) );
  OAI21_X1 U140 ( .B1(n872), .B2(n857), .A(n121), .ZN(n520) );
  BUF_X1 U141 ( .A(n3), .Z(n118) );
  INV_X1 U142 ( .A(n119), .ZN(n121) );
  NOR2_X1 U143 ( .A1(n453), .A2(n508), .ZN(n480) );
  AOI21_X1 U144 ( .B1(n480), .B2(N62), .A(n857), .ZN(n475) );
  OAI21_X1 U145 ( .B1(n518), .B2(n521), .A(n6), .ZN(N893) );
  OAI21_X1 U146 ( .B1(n518), .B2(n523), .A(n6), .ZN(N891) );
  OAI21_X1 U147 ( .B1(n518), .B2(n525), .A(n6), .ZN(N889) );
  OAI21_X1 U148 ( .B1(n518), .B2(n527), .A(n6), .ZN(N887) );
  OAI21_X1 U149 ( .B1(n518), .B2(n519), .A(n6), .ZN(N894) );
  OAI21_X1 U150 ( .B1(n518), .B2(n522), .A(n6), .ZN(N892) );
  OAI21_X1 U151 ( .B1(n518), .B2(n524), .A(n6), .ZN(N890) );
  OAI21_X1 U152 ( .B1(n518), .B2(n526), .A(n6), .ZN(N888) );
  OAI21_X1 U153 ( .B1(n521), .B2(n531), .A(n4), .ZN(N869) );
  OAI21_X1 U154 ( .B1(n523), .B2(n531), .A(n4), .ZN(N867) );
  OAI21_X1 U155 ( .B1(n525), .B2(n531), .A(n4), .ZN(N865) );
  OAI21_X1 U156 ( .B1(n527), .B2(n531), .A(n4), .ZN(N863) );
  OAI21_X1 U157 ( .B1(n519), .B2(n531), .A(n4), .ZN(N870) );
  OAI21_X1 U158 ( .B1(n522), .B2(n531), .A(n4), .ZN(N868) );
  OAI21_X1 U159 ( .B1(n524), .B2(n531), .A(n4), .ZN(N866) );
  OAI21_X1 U160 ( .B1(n526), .B2(n531), .A(n4), .ZN(N864) );
  OAI21_X1 U161 ( .B1(n521), .B2(n530), .A(n5), .ZN(N877) );
  OAI21_X1 U162 ( .B1(n521), .B2(n529), .A(n5), .ZN(N885) );
  OAI21_X1 U163 ( .B1(n523), .B2(n530), .A(n5), .ZN(N875) );
  OAI21_X1 U164 ( .B1(n523), .B2(n529), .A(n5), .ZN(N883) );
  OAI21_X1 U165 ( .B1(n525), .B2(n530), .A(n4), .ZN(N873) );
  OAI21_X1 U166 ( .B1(n525), .B2(n529), .A(n5), .ZN(N881) );
  OAI21_X1 U167 ( .B1(n527), .B2(n530), .A(n4), .ZN(N871) );
  OAI21_X1 U168 ( .B1(n527), .B2(n529), .A(n5), .ZN(N879) );
  OAI21_X1 U169 ( .B1(n519), .B2(n530), .A(n5), .ZN(N878) );
  OAI21_X1 U170 ( .B1(n519), .B2(n529), .A(n5), .ZN(N886) );
  OAI21_X1 U171 ( .B1(n522), .B2(n530), .A(n5), .ZN(N876) );
  OAI21_X1 U172 ( .B1(n522), .B2(n529), .A(n5), .ZN(N884) );
  OAI21_X1 U173 ( .B1(n524), .B2(n530), .A(n4), .ZN(N874) );
  OAI21_X1 U174 ( .B1(n524), .B2(n529), .A(n5), .ZN(N882) );
  OAI21_X1 U175 ( .B1(n526), .B2(n530), .A(n4), .ZN(N872) );
  OAI21_X1 U176 ( .B1(n526), .B2(n529), .A(n5), .ZN(N880) );
  INV_X1 U177 ( .A(N62), .ZN(n873) );
  BUF_X1 U178 ( .A(n1), .Z(n34) );
  BUF_X1 U179 ( .A(n1), .Z(n33) );
  INV_X1 U180 ( .A(n492), .ZN(n198) );
  INV_X1 U181 ( .A(n453), .ZN(n872) );
  BUF_X1 U182 ( .A(n282), .Z(n13) );
  BUF_X1 U183 ( .A(n280), .Z(n16) );
  BUF_X1 U184 ( .A(n282), .Z(n14) );
  BUF_X1 U185 ( .A(n280), .Z(n17) );
  BUF_X1 U186 ( .A(n286), .Z(n7) );
  BUF_X1 U187 ( .A(n284), .Z(n10) );
  BUF_X1 U188 ( .A(n286), .Z(n8) );
  BUF_X1 U189 ( .A(n284), .Z(n11) );
  INV_X1 U190 ( .A(n455), .ZN(n272) );
  INV_X1 U191 ( .A(n461), .ZN(n857) );
  BUF_X1 U192 ( .A(n282), .Z(n15) );
  BUF_X1 U193 ( .A(n280), .Z(n18) );
  BUF_X1 U194 ( .A(n286), .Z(n9) );
  BUF_X1 U195 ( .A(n284), .Z(n12) );
  BUF_X1 U196 ( .A(n1), .Z(n28) );
  BUF_X1 U197 ( .A(n1), .Z(n29) );
  BUF_X1 U198 ( .A(n1), .Z(n30) );
  BUF_X1 U199 ( .A(n1), .Z(n32) );
  BUF_X1 U200 ( .A(n1), .Z(n31) );
  BUF_X1 U201 ( .A(n1), .Z(n25) );
  BUF_X1 U202 ( .A(n1), .Z(n26) );
  BUF_X1 U203 ( .A(n1), .Z(n27) );
  BUF_X1 U204 ( .A(n1), .Z(n35) );
  BUF_X1 U205 ( .A(host_reset), .Z(n119) );
  BUF_X1 U206 ( .A(host_reset), .Z(n120) );
  INV_X1 U207 ( .A(n458), .ZN(n162) );
  AOI22_X1 U208 ( .A1(N257), .A2(n272), .B1(num_warps_out[4]), .B2(n455), .ZN(
        n458) );
  INV_X1 U209 ( .A(n456), .ZN(n170) );
  AOI22_X1 U210 ( .A1(N255), .A2(n272), .B1(num_warps_out[2]), .B2(n455), .ZN(
        n456) );
  INV_X1 U211 ( .A(n452), .ZN(n183) );
  AOI22_X1 U212 ( .A1(N91), .A2(n438), .B1(shmem_addr_i[13]), .B2(n439), .ZN(
        n452) );
  INV_X1 U213 ( .A(n454), .ZN(n174) );
  AOI22_X1 U214 ( .A1(N254), .A2(n272), .B1(num_warps_out[1]), .B2(n455), .ZN(
        n454) );
  INV_X1 U215 ( .A(n457), .ZN(n166) );
  AOI22_X1 U216 ( .A1(N256), .A2(n272), .B1(num_warps_out[3]), .B2(n455), .ZN(
        n457) );
  INV_X1 U217 ( .A(n468), .ZN(n168) );
  AOI22_X1 U218 ( .A1(n50), .A2(warp_pool_addr_out[3]), .B1(n32), .B2(
        warp_id_o[3]), .ZN(n468) );
  INV_X1 U219 ( .A(n463), .ZN(n169) );
  AOI22_X1 U220 ( .A1(n49), .A2(warp_state_addr_out[3]), .B1(n31), .B2(
        warp_id_o[3]), .ZN(n463) );
  INV_X1 U221 ( .A(n469), .ZN(n172) );
  AOI22_X1 U222 ( .A1(n50), .A2(warp_pool_addr_out[2]), .B1(n32), .B2(
        warp_id_o[2]), .ZN(n469) );
  INV_X1 U223 ( .A(n464), .ZN(n173) );
  AOI22_X1 U224 ( .A1(n49), .A2(warp_state_addr_out[2]), .B1(n31), .B2(
        warp_id_o[2]), .ZN(n464) );
  INV_X1 U225 ( .A(n470), .ZN(n176) );
  AOI22_X1 U226 ( .A1(n50), .A2(warp_pool_addr_out[1]), .B1(n32), .B2(
        warp_id_o[1]), .ZN(n470) );
  INV_X1 U227 ( .A(n465), .ZN(n177) );
  AOI22_X1 U228 ( .A1(n49), .A2(warp_state_addr_out[1]), .B1(n31), .B2(
        warp_id_o[1]), .ZN(n465) );
  INV_X1 U229 ( .A(n467), .ZN(n164) );
  AOI22_X1 U230 ( .A1(n50), .A2(warp_pool_addr_out[4]), .B1(n32), .B2(
        warp_id_o[4]), .ZN(n467) );
  INV_X1 U231 ( .A(n462), .ZN(n165) );
  AOI22_X1 U232 ( .A1(n48), .A2(warp_state_addr_out[4]), .B1(n30), .B2(
        warp_id_o[4]), .ZN(n462) );
  INV_X1 U233 ( .A(warps_per_block_in[4]), .ZN(n137) );
  INV_X1 U234 ( .A(n502), .ZN(n818) );
  AOI22_X1 U235 ( .A1(warps_per_block_cnt[4]), .A2(n496), .B1(n495), .B2(N96), 
        .ZN(n502) );
  INV_X1 U236 ( .A(n503), .ZN(n817) );
  AOI22_X1 U237 ( .A1(warps_per_block_cnt[3]), .A2(n496), .B1(n495), .B2(N95), 
        .ZN(n503) );
  INV_X1 U238 ( .A(n504), .ZN(n816) );
  AOI22_X1 U239 ( .A1(warps_per_block_cnt[2]), .A2(n496), .B1(n495), .B2(N94), 
        .ZN(n504) );
  INV_X1 U240 ( .A(n505), .ZN(n279) );
  AOI22_X1 U241 ( .A1(warps_per_block_cnt[1]), .A2(n496), .B1(n495), .B2(N93), 
        .ZN(n505) );
  INV_X1 U242 ( .A(n506), .ZN(n278) );
  AOI22_X1 U243 ( .A1(warps_per_block_cnt[0]), .A2(n496), .B1(n495), .B2(N92), 
        .ZN(n506) );
  NAND4_X1 U244 ( .A1(n455), .A2(n19), .A3(n511), .A4(n512), .ZN(n492) );
  AOI21_X1 U245 ( .B1(en), .B2(n857), .A(n413), .ZN(n512) );
  OAI21_X1 U246 ( .B1(n508), .B2(N62), .A(n872), .ZN(n511) );
  INV_X1 U247 ( .A(n130), .ZN(n138) );
  AOI21_X1 U248 ( .B1(n141), .B2(num_blocks_in[3]), .A(n874), .ZN(n508) );
  INV_X1 U249 ( .A(n513), .ZN(n874) );
  OAI222_X1 U250 ( .A1(n875), .A2(n142), .B1(num_blocks_in[2]), .B2(n514), 
        .C1(num_blocks_in[3]), .C2(n141), .ZN(n513) );
  INV_X1 U251 ( .A(n515), .ZN(n875) );
  OAI21_X1 U252 ( .B1(block_num_cnt[1]), .B2(n453), .A(n486), .ZN(n484) );
  AOI21_X1 U253 ( .B1(n145), .B2(n872), .A(n488), .ZN(n486) );
  OAI22_X1 U254 ( .A1(n155), .A2(n274), .B1(n473), .B2(n145), .ZN(n807) );
  OAI21_X1 U255 ( .B1(n516), .B2(num_blocks_in[1]), .A(n517), .ZN(n515) );
  OAI21_X1 U256 ( .B1(block_num_cnt[0]), .B2(n876), .A(block_num_cnt[1]), .ZN(
        n517) );
  NOR3_X1 U257 ( .A1(n876), .A2(block_num_cnt[1]), .A3(block_num_cnt[0]), .ZN(
        n516) );
  INV_X1 U258 ( .A(num_blocks_in[0]), .ZN(n876) );
  OAI22_X1 U259 ( .A1(n152), .A2(n274), .B1(n141), .B2(n473), .ZN(n801) );
  OAI22_X1 U260 ( .A1(n153), .A2(n274), .B1(n142), .B2(n473), .ZN(n800) );
  OAI22_X1 U261 ( .A1(n154), .A2(n274), .B1(n143), .B2(n473), .ZN(n799) );
  OAI22_X1 U262 ( .A1(n412), .A2(n175), .B1(n199), .B2(n270), .ZN(n725) );
  INV_X1 U263 ( .A(warp_id_o[1]), .ZN(n175) );
  OAI22_X1 U264 ( .A1(n412), .A2(n171), .B1(n199), .B2(n269), .ZN(n726) );
  INV_X1 U265 ( .A(warp_id_o[2]), .ZN(n171) );
  OAI22_X1 U266 ( .A1(n412), .A2(n167), .B1(n199), .B2(n268), .ZN(n727) );
  INV_X1 U267 ( .A(warp_id_o[3]), .ZN(n167) );
  OAI22_X1 U268 ( .A1(n412), .A2(n163), .B1(n199), .B2(n267), .ZN(n728) );
  INV_X1 U269 ( .A(warp_id_o[4]), .ZN(n163) );
  OAI22_X1 U270 ( .A1(n276), .A2(n142), .B1(n483), .B2(n485), .ZN(n809) );
  INV_X1 U271 ( .A(n484), .ZN(n276) );
  OAI22_X1 U272 ( .A1(n839), .A2(n21), .B1(N877), .B2(n220), .ZN(n581) );
  OAI22_X1 U273 ( .A1(n839), .A2(n21), .B1(N877), .B2(n252), .ZN(n549) );
  OAI22_X1 U274 ( .A1(n847), .A2(n19), .B1(N885), .B2(n212), .ZN(n573) );
  OAI22_X1 U275 ( .A1(n847), .A2(n22), .B1(N885), .B2(n244), .ZN(n541) );
  OAI22_X1 U276 ( .A1(n837), .A2(n21), .B1(N875), .B2(n222), .ZN(n583) );
  OAI22_X1 U277 ( .A1(n837), .A2(n19), .B1(N875), .B2(n254), .ZN(n551) );
  OAI22_X1 U278 ( .A1(n845), .A2(n20), .B1(N883), .B2(n214), .ZN(n575) );
  OAI22_X1 U279 ( .A1(n845), .A2(n20), .B1(N883), .B2(n246), .ZN(n543) );
  OAI22_X1 U280 ( .A1(n835), .A2(n21), .B1(N873), .B2(n224), .ZN(n585) );
  OAI22_X1 U281 ( .A1(n835), .A2(n19), .B1(N873), .B2(n256), .ZN(n553) );
  OAI22_X1 U282 ( .A1(n843), .A2(n21), .B1(N881), .B2(n216), .ZN(n577) );
  OAI22_X1 U283 ( .A1(n843), .A2(n21), .B1(N881), .B2(n248), .ZN(n545) );
  OAI22_X1 U284 ( .A1(n833), .A2(n22), .B1(N871), .B2(n226), .ZN(n587) );
  OAI22_X1 U285 ( .A1(n833), .A2(n19), .B1(N871), .B2(n258), .ZN(n555) );
  OAI22_X1 U286 ( .A1(n841), .A2(n21), .B1(N879), .B2(n218), .ZN(n579) );
  OAI22_X1 U287 ( .A1(n841), .A2(n22), .B1(N879), .B2(n250), .ZN(n547) );
  OAI22_X1 U288 ( .A1(n840), .A2(n21), .B1(N878), .B2(n219), .ZN(n580) );
  OAI22_X1 U289 ( .A1(n840), .A2(n24), .B1(N878), .B2(n251), .ZN(n548) );
  OAI22_X1 U290 ( .A1(n848), .A2(n19), .B1(N886), .B2(n211), .ZN(n572) );
  OAI22_X1 U291 ( .A1(n848), .A2(n20), .B1(N886), .B2(n243), .ZN(n540) );
  OAI22_X1 U292 ( .A1(n838), .A2(n21), .B1(N876), .B2(n221), .ZN(n582) );
  OAI22_X1 U293 ( .A1(n838), .A2(n19), .B1(N876), .B2(n253), .ZN(n550) );
  OAI22_X1 U294 ( .A1(n846), .A2(n20), .B1(N884), .B2(n213), .ZN(n574) );
  OAI22_X1 U295 ( .A1(n846), .A2(n24), .B1(N884), .B2(n245), .ZN(n542) );
  OAI22_X1 U296 ( .A1(n836), .A2(n21), .B1(N874), .B2(n223), .ZN(n584) );
  OAI22_X1 U297 ( .A1(n836), .A2(n19), .B1(N874), .B2(n255), .ZN(n552) );
  OAI22_X1 U298 ( .A1(n844), .A2(n21), .B1(N882), .B2(n215), .ZN(n576) );
  OAI22_X1 U299 ( .A1(n844), .A2(n23), .B1(N882), .B2(n247), .ZN(n544) );
  OAI22_X1 U300 ( .A1(n834), .A2(n20), .B1(N872), .B2(n225), .ZN(n586) );
  OAI22_X1 U301 ( .A1(n834), .A2(n19), .B1(N872), .B2(n257), .ZN(n554) );
  OAI22_X1 U302 ( .A1(n842), .A2(n21), .B1(N880), .B2(n217), .ZN(n578) );
  OAI22_X1 U303 ( .A1(n842), .A2(n19), .B1(N880), .B2(n249), .ZN(n546) );
  OAI22_X1 U304 ( .A1(n831), .A2(n22), .B1(N869), .B2(n228), .ZN(n589) );
  OAI22_X1 U305 ( .A1(n831), .A2(n19), .B1(N869), .B2(n260), .ZN(n557) );
  OAI22_X1 U306 ( .A1(n829), .A2(n20), .B1(N867), .B2(n230), .ZN(n591) );
  OAI22_X1 U307 ( .A1(n829), .A2(n20), .B1(N867), .B2(n262), .ZN(n559) );
  OAI22_X1 U308 ( .A1(n827), .A2(n21), .B1(N865), .B2(n232), .ZN(n593) );
  OAI22_X1 U309 ( .A1(n827), .A2(n20), .B1(N865), .B2(n264), .ZN(n561) );
  OAI22_X1 U310 ( .A1(n825), .A2(n21), .B1(N863), .B2(n234), .ZN(n595) );
  OAI22_X1 U311 ( .A1(n825), .A2(n20), .B1(N863), .B2(n266), .ZN(n563) );
  OAI22_X1 U312 ( .A1(n832), .A2(n22), .B1(N870), .B2(n227), .ZN(n588) );
  OAI22_X1 U314 ( .A1(n832), .A2(n19), .B1(N870), .B2(n259), .ZN(n556) );
  OAI22_X1 U315 ( .A1(n830), .A2(n20), .B1(N868), .B2(n229), .ZN(n590) );
  OAI22_X1 U316 ( .A1(n830), .A2(n19), .B1(N868), .B2(n261), .ZN(n558) );
  OAI22_X1 U317 ( .A1(n828), .A2(n24), .B1(N866), .B2(n231), .ZN(n592) );
  OAI22_X1 U318 ( .A1(n828), .A2(n20), .B1(N866), .B2(n263), .ZN(n560) );
  OAI22_X1 U319 ( .A1(n826), .A2(n23), .B1(N864), .B2(n233), .ZN(n594) );
  OAI22_X1 U320 ( .A1(n826), .A2(n20), .B1(N864), .B2(n265), .ZN(n562) );
  INV_X1 U321 ( .A(n428), .ZN(n140) );
  AOI22_X1 U322 ( .A1(gprs_base_addr_o[8]), .A2(n25), .B1(
        warp_pool_wr_data_out[105]), .B2(n39), .ZN(n428) );
  INV_X1 U323 ( .A(n431), .ZN(n157) );
  AOI22_X1 U324 ( .A1(gprs_base_addr_o[5]), .A2(n26), .B1(
        warp_pool_wr_data_out[102]), .B2(n39), .ZN(n431) );
  OAI22_X1 U325 ( .A1(n855), .A2(n20), .B1(N893), .B2(n204), .ZN(n565) );
  OAI22_X1 U326 ( .A1(n855), .A2(n24), .B1(N893), .B2(n236), .ZN(n533) );
  OAI22_X1 U327 ( .A1(n853), .A2(n20), .B1(N891), .B2(n206), .ZN(n567) );
  OAI22_X1 U328 ( .A1(n853), .A2(n21), .B1(N891), .B2(n238), .ZN(n535) );
  OAI22_X1 U329 ( .A1(n851), .A2(n21), .B1(N889), .B2(n208), .ZN(n569) );
  OAI22_X1 U330 ( .A1(n851), .A2(n20), .B1(N889), .B2(n240), .ZN(n537) );
  OAI22_X1 U331 ( .A1(n849), .A2(n21), .B1(N887), .B2(n210), .ZN(n571) );
  OAI22_X1 U332 ( .A1(n849), .A2(n22), .B1(N887), .B2(n242), .ZN(n539) );
  OAI22_X1 U333 ( .A1(n856), .A2(n20), .B1(N894), .B2(n203), .ZN(n564) );
  OAI22_X1 U334 ( .A1(n856), .A2(n19), .B1(N894), .B2(n235), .ZN(n532) );
  OAI22_X1 U335 ( .A1(n854), .A2(n20), .B1(N892), .B2(n205), .ZN(n566) );
  OAI22_X1 U336 ( .A1(n854), .A2(n23), .B1(N892), .B2(n237), .ZN(n534) );
  OAI22_X1 U337 ( .A1(n852), .A2(n21), .B1(N890), .B2(n207), .ZN(n568) );
  OAI22_X1 U338 ( .A1(n852), .A2(n21), .B1(N890), .B2(n239), .ZN(n536) );
  OAI22_X1 U339 ( .A1(n850), .A2(n19), .B1(N888), .B2(n209), .ZN(n570) );
  OAI22_X1 U340 ( .A1(n850), .A2(n20), .B1(N888), .B2(n241), .ZN(n538) );
  OAI22_X1 U341 ( .A1(n486), .A2(n143), .B1(block_num_cnt[1]), .B2(n483), .ZN(
        n811) );
  OAI22_X1 U342 ( .A1(n36), .A2(n40), .B1(n24), .B2(n152), .ZN(n729) );
  OAI22_X1 U343 ( .A1(n37), .A2(n41), .B1(n23), .B2(n153), .ZN(n730) );
  OAI22_X1 U344 ( .A1(n36), .A2(n42), .B1(n22), .B2(n154), .ZN(n731) );
  AND2_X1 U345 ( .A1(warps_per_block_in[0]), .A2(n151), .ZN(n129) );
  OAI22_X1 U346 ( .A1(n202), .A2(n492), .B1(n198), .B2(n510), .ZN(n815) );
  NOR2_X1 U347 ( .A1(n38), .A2(n413), .ZN(n510) );
  OAI22_X1 U348 ( .A1(n37), .A2(n43), .B1(n19), .B2(n155), .ZN(n732) );
  OAI21_X1 U349 ( .B1(n473), .B2(n147), .A(n479), .ZN(n806) );
  OAI21_X1 U350 ( .B1(n473), .B2(n148), .A(n478), .ZN(n805) );
  OAI21_X1 U351 ( .B1(n473), .B2(n149), .A(n477), .ZN(n804) );
  OAI21_X1 U352 ( .B1(n473), .B2(n150), .A(n476), .ZN(n803) );
  OAI21_X1 U353 ( .B1(n473), .B2(n151), .A(n474), .ZN(n802) );
  OAI21_X1 U354 ( .B1(n201), .B2(n492), .A(n493), .ZN(n814) );
  OAI21_X1 U355 ( .B1(n480), .B2(n413), .A(n492), .ZN(n493) );
  OAI21_X1 U356 ( .B1(n831), .B2(n7), .A(n387), .ZN(n699) );
  OAI21_X1 U357 ( .B1(n831), .B2(n10), .A(n386), .ZN(n698) );
  OAI21_X1 U358 ( .B1(n831), .B2(n13), .A(n385), .ZN(n697) );
  OAI21_X1 U359 ( .B1(n831), .B2(n16), .A(n384), .ZN(n696) );
  OAI21_X1 U360 ( .B1(n839), .B2(n8), .A(n355), .ZN(n667) );
  OAI21_X1 U361 ( .B1(n839), .B2(n11), .A(n354), .ZN(n666) );
  OAI21_X1 U362 ( .B1(n839), .B2(n14), .A(n353), .ZN(n665) );
  OAI21_X1 U363 ( .B1(n839), .B2(n17), .A(n352), .ZN(n664) );
  OAI21_X1 U364 ( .B1(n847), .B2(n8), .A(n323), .ZN(n635) );
  OAI21_X1 U365 ( .B1(n847), .B2(n11), .A(n322), .ZN(n634) );
  OAI21_X1 U366 ( .B1(n847), .B2(n14), .A(n321), .ZN(n633) );
  OAI21_X1 U367 ( .B1(n847), .B2(n17), .A(n320), .ZN(n632) );
  OAI21_X1 U368 ( .B1(n829), .B2(n7), .A(n395), .ZN(n707) );
  OAI21_X1 U369 ( .B1(n829), .B2(n10), .A(n394), .ZN(n706) );
  OAI21_X1 U370 ( .B1(n829), .B2(n13), .A(n393), .ZN(n705) );
  OAI21_X1 U371 ( .B1(n829), .B2(n16), .A(n392), .ZN(n704) );
  OAI21_X1 U372 ( .B1(n837), .B2(n8), .A(n363), .ZN(n675) );
  OAI21_X1 U373 ( .B1(n837), .B2(n11), .A(n362), .ZN(n674) );
  OAI21_X1 U374 ( .B1(n837), .B2(n14), .A(n361), .ZN(n673) );
  OAI21_X1 U375 ( .B1(n837), .B2(n17), .A(n360), .ZN(n672) );
  OAI21_X1 U376 ( .B1(n845), .B2(n8), .A(n331), .ZN(n643) );
  OAI21_X1 U377 ( .B1(n845), .B2(n11), .A(n330), .ZN(n642) );
  OAI21_X1 U378 ( .B1(n845), .B2(n14), .A(n329), .ZN(n641) );
  OAI21_X1 U379 ( .B1(n845), .B2(n17), .A(n328), .ZN(n640) );
  OAI21_X1 U380 ( .B1(n827), .B2(n7), .A(n403), .ZN(n715) );
  OAI21_X1 U381 ( .B1(n827), .B2(n10), .A(n402), .ZN(n714) );
  OAI21_X1 U382 ( .B1(n827), .B2(n13), .A(n401), .ZN(n713) );
  OAI21_X1 U383 ( .B1(n827), .B2(n16), .A(n400), .ZN(n712) );
  OAI21_X1 U384 ( .B1(n835), .B2(n7), .A(n371), .ZN(n683) );
  OAI21_X1 U385 ( .B1(n835), .B2(n10), .A(n370), .ZN(n682) );
  OAI21_X1 U386 ( .B1(n835), .B2(n13), .A(n369), .ZN(n681) );
  OAI21_X1 U387 ( .B1(n835), .B2(n16), .A(n368), .ZN(n680) );
  OAI21_X1 U388 ( .B1(n843), .B2(n8), .A(n339), .ZN(n651) );
  OAI21_X1 U389 ( .B1(n843), .B2(n11), .A(n338), .ZN(n650) );
  OAI21_X1 U390 ( .B1(n843), .B2(n14), .A(n337), .ZN(n649) );
  OAI21_X1 U391 ( .B1(n843), .B2(n17), .A(n336), .ZN(n648) );
  OAI21_X1 U392 ( .B1(n825), .B2(n7), .A(n411), .ZN(n723) );
  OAI21_X1 U393 ( .B1(n825), .B2(n10), .A(n410), .ZN(n722) );
  OAI21_X1 U394 ( .B1(n825), .B2(n13), .A(n409), .ZN(n721) );
  OAI21_X1 U395 ( .B1(n825), .B2(n16), .A(n408), .ZN(n720) );
  OAI21_X1 U396 ( .B1(n833), .B2(n7), .A(n379), .ZN(n691) );
  OAI21_X1 U397 ( .B1(n833), .B2(n10), .A(n378), .ZN(n690) );
  OAI21_X1 U398 ( .B1(n833), .B2(n13), .A(n377), .ZN(n689) );
  OAI21_X1 U399 ( .B1(n833), .B2(n16), .A(n376), .ZN(n688) );
  OAI21_X1 U400 ( .B1(n841), .B2(n8), .A(n347), .ZN(n659) );
  OAI21_X1 U401 ( .B1(n841), .B2(n11), .A(n346), .ZN(n658) );
  OAI21_X1 U402 ( .B1(n841), .B2(n14), .A(n345), .ZN(n657) );
  OAI21_X1 U403 ( .B1(n841), .B2(n17), .A(n344), .ZN(n656) );
  OAI21_X1 U404 ( .B1(n832), .B2(n7), .A(n383), .ZN(n695) );
  OAI21_X1 U405 ( .B1(n832), .B2(n10), .A(n382), .ZN(n694) );
  OAI21_X1 U406 ( .B1(n832), .B2(n13), .A(n381), .ZN(n693) );
  OAI21_X1 U407 ( .B1(n832), .B2(n16), .A(n380), .ZN(n692) );
  OAI21_X1 U408 ( .B1(n840), .B2(n8), .A(n351), .ZN(n663) );
  OAI21_X1 U409 ( .B1(n840), .B2(n11), .A(n350), .ZN(n662) );
  OAI21_X1 U410 ( .B1(n840), .B2(n14), .A(n349), .ZN(n661) );
  OAI21_X1 U411 ( .B1(n840), .B2(n17), .A(n348), .ZN(n660) );
  OAI21_X1 U412 ( .B1(n848), .B2(n8), .A(n319), .ZN(n631) );
  OAI21_X1 U413 ( .B1(n848), .B2(n11), .A(n318), .ZN(n630) );
  OAI21_X1 U414 ( .B1(n848), .B2(n14), .A(n317), .ZN(n629) );
  OAI21_X1 U415 ( .B1(n848), .B2(n17), .A(n316), .ZN(n628) );
  OAI21_X1 U416 ( .B1(n830), .B2(n7), .A(n391), .ZN(n703) );
  OAI21_X1 U417 ( .B1(n830), .B2(n10), .A(n390), .ZN(n702) );
  OAI21_X1 U418 ( .B1(n830), .B2(n13), .A(n389), .ZN(n701) );
  OAI21_X1 U419 ( .B1(n830), .B2(n16), .A(n388), .ZN(n700) );
  OAI21_X1 U420 ( .B1(n838), .B2(n8), .A(n359), .ZN(n671) );
  OAI21_X1 U421 ( .B1(n838), .B2(n11), .A(n358), .ZN(n670) );
  OAI21_X1 U422 ( .B1(n838), .B2(n14), .A(n357), .ZN(n669) );
  OAI21_X1 U423 ( .B1(n838), .B2(n17), .A(n356), .ZN(n668) );
  OAI21_X1 U424 ( .B1(n846), .B2(n8), .A(n327), .ZN(n639) );
  OAI21_X1 U425 ( .B1(n846), .B2(n11), .A(n326), .ZN(n638) );
  OAI21_X1 U426 ( .B1(n846), .B2(n14), .A(n325), .ZN(n637) );
  OAI21_X1 U427 ( .B1(n846), .B2(n17), .A(n324), .ZN(n636) );
  OAI21_X1 U428 ( .B1(n828), .B2(n7), .A(n399), .ZN(n711) );
  OAI21_X1 U430 ( .B1(n828), .B2(n10), .A(n398), .ZN(n710) );
  OAI21_X1 U431 ( .B1(n828), .B2(n13), .A(n397), .ZN(n709) );
  OAI21_X1 U432 ( .B1(n828), .B2(n16), .A(n396), .ZN(n708) );
  OAI21_X1 U433 ( .B1(n836), .B2(n7), .A(n367), .ZN(n679) );
  OAI21_X1 U434 ( .B1(n836), .B2(n10), .A(n366), .ZN(n678) );
  OAI21_X1 U435 ( .B1(n836), .B2(n13), .A(n365), .ZN(n677) );
  OAI21_X1 U436 ( .B1(n836), .B2(n16), .A(n364), .ZN(n676) );
  OAI21_X1 U437 ( .B1(n844), .B2(n8), .A(n335), .ZN(n647) );
  OAI21_X1 U438 ( .B1(n844), .B2(n11), .A(n334), .ZN(n646) );
  OAI21_X1 U439 ( .B1(n844), .B2(n14), .A(n333), .ZN(n645) );
  OAI21_X1 U440 ( .B1(n844), .B2(n17), .A(n332), .ZN(n644) );
  OAI21_X1 U441 ( .B1(n826), .B2(n7), .A(n407), .ZN(n719) );
  OAI21_X1 U442 ( .B1(n826), .B2(n10), .A(n406), .ZN(n718) );
  OAI21_X1 U443 ( .B1(n826), .B2(n13), .A(n405), .ZN(n717) );
  OAI21_X1 U444 ( .B1(n826), .B2(n16), .A(n404), .ZN(n716) );
  OAI21_X1 U445 ( .B1(n834), .B2(n7), .A(n375), .ZN(n687) );
  OAI21_X1 U446 ( .B1(n834), .B2(n10), .A(n374), .ZN(n686) );
  OAI21_X1 U447 ( .B1(n834), .B2(n13), .A(n373), .ZN(n685) );
  OAI21_X1 U448 ( .B1(n834), .B2(n16), .A(n372), .ZN(n684) );
  OAI21_X1 U449 ( .B1(n842), .B2(n8), .A(n343), .ZN(n655) );
  OAI21_X1 U450 ( .B1(n842), .B2(n11), .A(n342), .ZN(n654) );
  OAI21_X1 U451 ( .B1(n842), .B2(n14), .A(n341), .ZN(n653) );
  OAI21_X1 U452 ( .B1(n842), .B2(n17), .A(n340), .ZN(n652) );
  OAI21_X1 U453 ( .B1(n38), .B2(n90), .A(n23), .ZN(n771) );
  OAI21_X1 U454 ( .B1(n37), .B2(n78), .A(n23), .ZN(n759) );
  OAI21_X1 U455 ( .B1(n37), .B2(n75), .A(n23), .ZN(n756) );
  OAI21_X1 U456 ( .B1(n37), .B2(n74), .A(n23), .ZN(n755) );
  OAI21_X1 U457 ( .B1(n37), .B2(n73), .A(n23), .ZN(n754) );
  OAI21_X1 U458 ( .B1(n37), .B2(n72), .A(n23), .ZN(n753) );
  OAI21_X1 U459 ( .B1(n36), .B2(n71), .A(n23), .ZN(n752) );
  OAI21_X1 U460 ( .B1(n36), .B2(n70), .A(n23), .ZN(n751) );
  OAI21_X1 U461 ( .B1(n36), .B2(n69), .A(n23), .ZN(n750) );
  OAI21_X1 U462 ( .B1(n36), .B2(n67), .A(n23), .ZN(n748) );
  OAI21_X1 U463 ( .B1(n36), .B2(n115), .A(n20), .ZN(n796) );
  OAI21_X1 U464 ( .B1(n37), .B2(n57), .A(n22), .ZN(n738) );
  OAI21_X1 U465 ( .B1(n36), .B2(n56), .A(n22), .ZN(n737) );
  OAI21_X1 U466 ( .B1(n37), .B2(n55), .A(n20), .ZN(n736) );
  OAI21_X1 U467 ( .B1(n36), .B2(n54), .A(n23), .ZN(n735) );
  OAI21_X1 U468 ( .B1(n37), .B2(n53), .A(n24), .ZN(n734) );
  OAI21_X1 U469 ( .B1(n36), .B2(n116), .A(n23), .ZN(n733) );
  NOR2_X1 U470 ( .A1(block_num_cnt[2]), .A2(n515), .ZN(n514) );
  OAI21_X1 U471 ( .B1(n36), .B2(n109), .A(n21), .ZN(n790) );
  OAI21_X1 U472 ( .B1(n37), .B2(n108), .A(n21), .ZN(n789) );
  OAI21_X1 U473 ( .B1(n36), .B2(n107), .A(n22), .ZN(n788) );
  OAI21_X1 U474 ( .B1(n37), .B2(n106), .A(n24), .ZN(n787) );
  OAI21_X1 U475 ( .B1(n36), .B2(n105), .A(n23), .ZN(n786) );
  OAI21_X1 U476 ( .B1(n37), .B2(n104), .A(n19), .ZN(n785) );
  OAI21_X1 U477 ( .B1(n36), .B2(n103), .A(n19), .ZN(n784) );
  OAI21_X1 U478 ( .B1(n38), .B2(n102), .A(n21), .ZN(n783) );
  OAI21_X1 U479 ( .B1(n38), .B2(n101), .A(n24), .ZN(n782) );
  OAI21_X1 U480 ( .B1(n38), .B2(n100), .A(n23), .ZN(n781) );
  OAI21_X1 U481 ( .B1(n38), .B2(n99), .A(n19), .ZN(n780) );
  OAI21_X1 U482 ( .B1(n38), .B2(n98), .A(n19), .ZN(n779) );
  OAI21_X1 U483 ( .B1(n38), .B2(n97), .A(n19), .ZN(n778) );
  OAI21_X1 U484 ( .B1(n38), .B2(n96), .A(n19), .ZN(n777) );
  OAI21_X1 U485 ( .B1(n38), .B2(n95), .A(n19), .ZN(n776) );
  OAI21_X1 U486 ( .B1(n38), .B2(n94), .A(n23), .ZN(n775) );
  OAI21_X1 U487 ( .B1(n38), .B2(n93), .A(n23), .ZN(n774) );
  OAI21_X1 U488 ( .B1(n38), .B2(n92), .A(n24), .ZN(n773) );
  OAI21_X1 U489 ( .B1(n38), .B2(n91), .A(n23), .ZN(n772) );
  OAI21_X1 U490 ( .B1(n38), .B2(n89), .A(n24), .ZN(n770) );
  OAI21_X1 U491 ( .B1(n38), .B2(n88), .A(n24), .ZN(n769) );
  OAI21_X1 U492 ( .B1(n38), .B2(n87), .A(n24), .ZN(n768) );
  OAI21_X1 U493 ( .B1(n38), .B2(n86), .A(n24), .ZN(n767) );
  OAI21_X1 U494 ( .B1(n38), .B2(n85), .A(n24), .ZN(n766) );
  OAI21_X1 U495 ( .B1(n38), .B2(n84), .A(n24), .ZN(n765) );
  OAI21_X1 U496 ( .B1(n37), .B2(n83), .A(n21), .ZN(n764) );
  OAI21_X1 U497 ( .B1(n37), .B2(n82), .A(n24), .ZN(n763) );
  OAI21_X1 U498 ( .B1(n37), .B2(n81), .A(n24), .ZN(n762) );
  OAI21_X1 U499 ( .B1(n37), .B2(n80), .A(n24), .ZN(n761) );
  OAI21_X1 U500 ( .B1(n37), .B2(n79), .A(n24), .ZN(n760) );
  OAI21_X1 U501 ( .B1(n37), .B2(n77), .A(n24), .ZN(n758) );
  OAI21_X1 U502 ( .B1(n37), .B2(n76), .A(n22), .ZN(n757) );
  OAI21_X1 U503 ( .B1(n36), .B2(n68), .A(n22), .ZN(n749) );
  OAI21_X1 U504 ( .B1(n36), .B2(n66), .A(n22), .ZN(n747) );
  OAI21_X1 U505 ( .B1(n36), .B2(n65), .A(n22), .ZN(n746) );
  OAI21_X1 U506 ( .B1(n37), .B2(n64), .A(n22), .ZN(n745) );
  OAI21_X1 U507 ( .B1(n36), .B2(n63), .A(n22), .ZN(n744) );
  OAI21_X1 U508 ( .B1(n36), .B2(n62), .A(n22), .ZN(n743) );
  OAI21_X1 U509 ( .B1(n36), .B2(n61), .A(n22), .ZN(n742) );
  OAI21_X1 U510 ( .B1(n36), .B2(n60), .A(n22), .ZN(n741) );
  OAI21_X1 U511 ( .B1(n36), .B2(n59), .A(n22), .ZN(n740) );
  OAI21_X1 U512 ( .B1(n36), .B2(n58), .A(n20), .ZN(n739) );
  OAI21_X1 U513 ( .B1(n855), .B2(n9), .A(n291), .ZN(n603) );
  OAI21_X1 U514 ( .B1(n855), .B2(n12), .A(n290), .ZN(n602) );
  OAI21_X1 U515 ( .B1(n855), .B2(n15), .A(n289), .ZN(n601) );
  OAI21_X1 U516 ( .B1(n855), .B2(n18), .A(n288), .ZN(n600) );
  OAI21_X1 U517 ( .B1(n853), .B2(n9), .A(n299), .ZN(n611) );
  OAI21_X1 U518 ( .B1(n853), .B2(n12), .A(n298), .ZN(n610) );
  OAI21_X1 U519 ( .B1(n853), .B2(n15), .A(n297), .ZN(n609) );
  OAI21_X1 U520 ( .B1(n853), .B2(n18), .A(n296), .ZN(n608) );
  OAI21_X1 U521 ( .B1(n851), .B2(n9), .A(n307), .ZN(n619) );
  OAI21_X1 U522 ( .B1(n851), .B2(n12), .A(n306), .ZN(n618) );
  OAI21_X1 U523 ( .B1(n851), .B2(n15), .A(n305), .ZN(n617) );
  OAI21_X1 U524 ( .B1(n851), .B2(n18), .A(n304), .ZN(n616) );
  OAI21_X1 U525 ( .B1(n849), .B2(n9), .A(n315), .ZN(n627) );
  OAI21_X1 U526 ( .B1(n849), .B2(n12), .A(n314), .ZN(n626) );
  OAI21_X1 U527 ( .B1(n849), .B2(n15), .A(n313), .ZN(n625) );
  OAI21_X1 U528 ( .B1(n849), .B2(n18), .A(n312), .ZN(n624) );
  OAI21_X1 U529 ( .B1(n856), .B2(n9), .A(n287), .ZN(n599) );
  OAI21_X1 U530 ( .B1(n856), .B2(n12), .A(n285), .ZN(n598) );
  OAI21_X1 U531 ( .B1(n856), .B2(n15), .A(n283), .ZN(n597) );
  OAI21_X1 U532 ( .B1(n856), .B2(n18), .A(n281), .ZN(n596) );
  OAI21_X1 U533 ( .B1(n854), .B2(n9), .A(n295), .ZN(n607) );
  OAI21_X1 U534 ( .B1(n854), .B2(n12), .A(n294), .ZN(n606) );
  OAI21_X1 U535 ( .B1(n854), .B2(n15), .A(n293), .ZN(n605) );
  OAI21_X1 U536 ( .B1(n854), .B2(n18), .A(n292), .ZN(n604) );
  OAI21_X1 U537 ( .B1(n852), .B2(n9), .A(n303), .ZN(n615) );
  OAI21_X1 U538 ( .B1(n852), .B2(n12), .A(n302), .ZN(n614) );
  OAI21_X1 U539 ( .B1(n852), .B2(n15), .A(n301), .ZN(n613) );
  OAI21_X1 U540 ( .B1(n852), .B2(n18), .A(n300), .ZN(n612) );
  OAI21_X1 U541 ( .B1(n850), .B2(n9), .A(n311), .ZN(n623) );
  OAI21_X1 U542 ( .B1(n850), .B2(n12), .A(n310), .ZN(n622) );
  OAI21_X1 U543 ( .B1(n850), .B2(n15), .A(n309), .ZN(n621) );
  OAI21_X1 U544 ( .B1(n850), .B2(n18), .A(n308), .ZN(n620) );
  OAI21_X1 U545 ( .B1(n145), .B2(n275), .A(n487), .ZN(n810) );
  OAI21_X1 U546 ( .B1(n481), .B2(n141), .A(n482), .ZN(n808) );
  NOR2_X1 U547 ( .A1(n872), .A2(n484), .ZN(n481) );
  OR3_X1 U548 ( .A1(n142), .A2(n143), .A3(n483), .ZN(n482) );
  INV_X1 U549 ( .A(warps_per_block_in[3]), .ZN(n136) );
  INV_X1 U550 ( .A(n494), .ZN(n824) );
  AOI22_X1 U551 ( .A1(N102), .A2(n495), .B1(warps_per_block_cnt[10]), .B2(n496), .ZN(n494) );
  INV_X1 U552 ( .A(n497), .ZN(n823) );
  AOI22_X1 U553 ( .A1(N101), .A2(n495), .B1(warps_per_block_cnt[9]), .B2(n496), 
        .ZN(n497) );
  INV_X1 U554 ( .A(n498), .ZN(n822) );
  AOI22_X1 U555 ( .A1(N100), .A2(n495), .B1(warps_per_block_cnt[8]), .B2(n496), 
        .ZN(n498) );
  INV_X1 U556 ( .A(n499), .ZN(n821) );
  AOI22_X1 U557 ( .A1(N99), .A2(n495), .B1(warps_per_block_cnt[7]), .B2(n496), 
        .ZN(n499) );
  INV_X1 U558 ( .A(n500), .ZN(n820) );
  AOI22_X1 U559 ( .A1(N98), .A2(n495), .B1(warps_per_block_cnt[6]), .B2(n496), 
        .ZN(n500) );
  INV_X1 U560 ( .A(n501), .ZN(n819) );
  AOI22_X1 U561 ( .A1(N97), .A2(n495), .B1(warps_per_block_cnt[5]), .B2(n496), 
        .ZN(n501) );
  INV_X1 U562 ( .A(n507), .ZN(n277) );
  AOI22_X1 U563 ( .A1(N103), .A2(n495), .B1(warps_per_block_cnt[11]), .B2(n496), .ZN(n507) );
  OAI22_X1 U564 ( .A1(n472), .A2(n453), .B1(n273), .B2(n156), .ZN(n798) );
  INV_X1 U565 ( .A(n472), .ZN(n273) );
  NOR2_X1 U566 ( .A1(n274), .A2(n413), .ZN(n472) );
  INV_X1 U567 ( .A(n437), .ZN(n196) );
  AOI22_X1 U568 ( .A1(N78), .A2(n438), .B1(shmem_addr_i[0]), .B2(n439), .ZN(
        n437) );
  INV_X1 U569 ( .A(n440), .ZN(n195) );
  AOI22_X1 U570 ( .A1(N79), .A2(n438), .B1(shmem_addr_i[1]), .B2(n439), .ZN(
        n440) );
  INV_X1 U571 ( .A(n441), .ZN(n194) );
  AOI22_X1 U572 ( .A1(N80), .A2(n438), .B1(shmem_addr_i[2]), .B2(n439), .ZN(
        n441) );
  INV_X1 U573 ( .A(n442), .ZN(n193) );
  AOI22_X1 U574 ( .A1(N81), .A2(n438), .B1(shmem_addr_i[3]), .B2(n439), .ZN(
        n442) );
  INV_X1 U575 ( .A(n443), .ZN(n192) );
  AOI22_X1 U576 ( .A1(N82), .A2(n438), .B1(shmem_addr_i[4]), .B2(n439), .ZN(
        n443) );
  INV_X1 U577 ( .A(n444), .ZN(n191) );
  AOI22_X1 U578 ( .A1(N83), .A2(n438), .B1(shmem_addr_i[5]), .B2(n439), .ZN(
        n444) );
  INV_X1 U579 ( .A(n445), .ZN(n190) );
  AOI22_X1 U580 ( .A1(N84), .A2(n438), .B1(shmem_addr_i[6]), .B2(n439), .ZN(
        n445) );
  INV_X1 U581 ( .A(n446), .ZN(n189) );
  AOI22_X1 U582 ( .A1(N85), .A2(n438), .B1(shmem_addr_i[7]), .B2(n439), .ZN(
        n446) );
  INV_X1 U583 ( .A(n447), .ZN(n188) );
  AOI22_X1 U584 ( .A1(N86), .A2(n438), .B1(shmem_addr_i[8]), .B2(n439), .ZN(
        n447) );
  INV_X1 U585 ( .A(n448), .ZN(n187) );
  AOI22_X1 U586 ( .A1(N87), .A2(n438), .B1(shmem_addr_i[9]), .B2(n439), .ZN(
        n448) );
  INV_X1 U587 ( .A(n449), .ZN(n186) );
  AOI22_X1 U588 ( .A1(N88), .A2(n438), .B1(shmem_addr_i[10]), .B2(n439), .ZN(
        n449) );
  INV_X1 U589 ( .A(n450), .ZN(n185) );
  AOI22_X1 U590 ( .A1(N89), .A2(n438), .B1(shmem_addr_i[11]), .B2(n439), .ZN(
        n450) );
  INV_X1 U591 ( .A(n451), .ZN(n184) );
  AOI22_X1 U592 ( .A1(N90), .A2(n438), .B1(shmem_addr_i[12]), .B2(n439), .ZN(
        n451) );
  INV_X1 U593 ( .A(n509), .ZN(n197) );
  AOI22_X1 U594 ( .A1(warp_generator_state_machine[2]), .A2(n198), .B1(n872), 
        .B2(n508), .ZN(n509) );
  INV_X1 U595 ( .A(n429), .ZN(n144) );
  AOI22_X1 U596 ( .A1(gprs_base_addr_o[7]), .A2(n25), .B1(
        warp_pool_wr_data_out[104]), .B2(n39), .ZN(n429) );
  INV_X1 U729 ( .A(n430), .ZN(n146) );
  AOI22_X1 U730 ( .A1(gprs_base_addr_o[6]), .A2(n25), .B1(
        warp_pool_wr_data_out[103]), .B2(n44), .ZN(n430) );
  INV_X1 U760 ( .A(n432), .ZN(n158) );
  AOI22_X1 U761 ( .A1(gprs_base_addr_o[4]), .A2(n26), .B1(
        warp_pool_wr_data_out[101]), .B2(n45), .ZN(n432) );
  INV_X1 U763 ( .A(n433), .ZN(n159) );
  AOI22_X1 U764 ( .A1(gprs_base_addr_o[3]), .A2(n25), .B1(
        warp_pool_wr_data_out[100]), .B2(n44), .ZN(n433) );
  INV_X1 U765 ( .A(n434), .ZN(n160) );
  AOI22_X1 U766 ( .A1(gprs_base_addr_o[2]), .A2(n26), .B1(
        warp_pool_wr_data_out[99]), .B2(n44), .ZN(n434) );
  OAI22_X1 U767 ( .A1(n412), .A2(n180), .B1(n199), .B2(n271), .ZN(n724) );
  INV_X1 U768 ( .A(warp_id_o[0]), .ZN(n180) );
  INV_X1 U769 ( .A(n436), .ZN(n178) );
  AOI22_X1 U770 ( .A1(gprs_base_addr_o[0]), .A2(n27), .B1(
        warp_pool_wr_data_out[97]), .B2(n44), .ZN(n436) );
  INV_X1 U771 ( .A(n435), .ZN(n161) );
  AOI22_X1 U772 ( .A1(gprs_base_addr_o[1]), .A2(n26), .B1(
        warp_pool_wr_data_out[98]), .B2(n39), .ZN(n435) );
  OAI21_X1 U773 ( .B1(n37), .B2(n114), .A(n22), .ZN(n795) );
  OAI21_X1 U774 ( .B1(n36), .B2(n113), .A(n20), .ZN(n794) );
  OAI21_X1 U775 ( .B1(n37), .B2(n112), .A(n24), .ZN(n793) );
  OAI21_X1 U776 ( .B1(n38), .B2(n111), .A(n23), .ZN(n792) );
  OAI21_X1 U777 ( .B1(n37), .B2(n110), .A(n20), .ZN(n791) );
  INV_X1 U778 ( .A(n459), .ZN(n179) );
  AOI22_X1 U779 ( .A1(n180), .A2(n272), .B1(num_warps_out[0]), .B2(n455), .ZN(
        n459) );
  INV_X1 U780 ( .A(n471), .ZN(n181) );
  AOI22_X1 U781 ( .A1(n51), .A2(warp_pool_addr_out[0]), .B1(n33), .B2(
        warp_id_o[0]), .ZN(n471) );
  INV_X1 U782 ( .A(n466), .ZN(n182) );
  AOI22_X1 U783 ( .A1(n49), .A2(warp_state_addr_out[0]), .B1(n31), .B2(
        warp_id_o[0]), .ZN(n466) );
  INV_X1 U784 ( .A(n427), .ZN(n871) );
  AOI22_X1 U785 ( .A1(n48), .A2(warp_pool_wr_data_out[110]), .B1(n29), .B2(
        shmem_addr_i[0]), .ZN(n427) );
  INV_X1 U786 ( .A(n426), .ZN(n870) );
  AOI22_X1 U787 ( .A1(n47), .A2(warp_pool_wr_data_out[111]), .B1(n29), .B2(
        shmem_addr_i[1]), .ZN(n426) );
  INV_X1 U788 ( .A(n425), .ZN(n869) );
  AOI22_X1 U789 ( .A1(n47), .A2(warp_pool_wr_data_out[112]), .B1(n30), .B2(
        shmem_addr_i[2]), .ZN(n425) );
  INV_X1 U790 ( .A(n424), .ZN(n868) );
  AOI22_X1 U791 ( .A1(n48), .A2(warp_pool_wr_data_out[113]), .B1(n29), .B2(
        shmem_addr_i[3]), .ZN(n424) );
  INV_X1 U792 ( .A(n423), .ZN(n867) );
  AOI22_X1 U793 ( .A1(n46), .A2(warp_pool_wr_data_out[114]), .B1(n28), .B2(
        shmem_addr_i[4]), .ZN(n423) );
  INV_X1 U794 ( .A(n422), .ZN(n866) );
  AOI22_X1 U795 ( .A1(n46), .A2(warp_pool_wr_data_out[115]), .B1(n30), .B2(
        shmem_addr_i[5]), .ZN(n422) );
  INV_X1 U796 ( .A(n421), .ZN(n865) );
  AOI22_X1 U797 ( .A1(n46), .A2(warp_pool_wr_data_out[116]), .B1(n28), .B2(
        shmem_addr_i[6]), .ZN(n421) );
  INV_X1 U798 ( .A(n420), .ZN(n864) );
  AOI22_X1 U799 ( .A1(n47), .A2(warp_pool_wr_data_out[117]), .B1(n30), .B2(
        shmem_addr_i[7]), .ZN(n420) );
  INV_X1 U800 ( .A(n419), .ZN(n863) );
  AOI22_X1 U801 ( .A1(n45), .A2(warp_pool_wr_data_out[118]), .B1(n28), .B2(
        shmem_addr_i[8]), .ZN(n419) );
  INV_X1 U802 ( .A(n418), .ZN(n862) );
  AOI22_X1 U803 ( .A1(n47), .A2(warp_pool_wr_data_out[119]), .B1(n28), .B2(
        shmem_addr_i[9]), .ZN(n418) );
  INV_X1 U804 ( .A(n417), .ZN(n861) );
  AOI22_X1 U805 ( .A1(n45), .A2(warp_pool_wr_data_out[120]), .B1(n27), .B2(
        shmem_addr_i[10]), .ZN(n417) );
  INV_X1 U806 ( .A(n416), .ZN(n860) );
  AOI22_X1 U807 ( .A1(n46), .A2(warp_pool_wr_data_out[121]), .B1(n29), .B2(
        shmem_addr_i[11]), .ZN(n416) );
  INV_X1 U808 ( .A(n415), .ZN(n859) );
  AOI22_X1 U809 ( .A1(n45), .A2(warp_pool_wr_data_out[122]), .B1(n27), .B2(
        shmem_addr_i[12]), .ZN(n415) );
  INV_X1 U810 ( .A(n414), .ZN(n858) );
  AOI22_X1 U811 ( .A1(n48), .A2(warp_pool_wr_data_out[123]), .B1(n27), .B2(
        shmem_addr_i[13]), .ZN(n414) );
  INV_X1 U812 ( .A(n34), .ZN(n23) );
  INV_X1 U813 ( .A(n119), .ZN(n122) );
  INV_X1 U814 ( .A(n119), .ZN(n123) );
  INV_X1 U815 ( .A(n119), .ZN(n124) );
  INV_X1 U816 ( .A(n119), .ZN(n125) );
  INV_X1 U817 ( .A(n120), .ZN(n126) );
  INV_X1 U818 ( .A(n120), .ZN(n127) );
  XOR2_X1 U819 ( .A(\add_155/carry[4] ), .B(warp_id_o[4]), .Z(N257) );
  OR4_X1 U820 ( .A1(warps_per_block_cnt[7]), .A2(warps_per_block_cnt[6]), .A3(
        warps_per_block_cnt[9]), .A4(warps_per_block_cnt[8]), .ZN(n135) );
  AND2_X1 U821 ( .A1(n150), .A2(n129), .ZN(n128) );
  OAI222_X1 U822 ( .A1(n129), .A2(n150), .B1(warps_per_block_in[1]), .B2(n128), 
        .C1(warps_per_block_in[2]), .C2(n149), .ZN(n130) );
  AOI221_X1 U823 ( .B1(n149), .B2(warps_per_block_in[2]), .C1(n148), .C2(
        warps_per_block_in[3]), .A(n138), .ZN(n131) );
  AOI221_X1 U824 ( .B1(n136), .B2(warps_per_block_cnt[3]), .C1(n137), .C2(
        warps_per_block_cnt[4]), .A(n131), .ZN(n132) );
  AOI221_X1 U825 ( .B1(n147), .B2(warps_per_block_in[4]), .C1(n2), .C2(
        warps_per_block_in[5]), .A(n132), .ZN(n133) );
  OAI21_X1 U826 ( .B1(warps_per_block_in[5]), .B2(n2), .A(n139), .ZN(n134) );
  NOR4_X1 U827 ( .A1(n135), .A2(n134), .A3(warps_per_block_cnt[11]), .A4(
        warps_per_block_cnt[10]), .ZN(N62) );
  NAND2_X1 U828 ( .A1(n413), .A2(n126), .ZN(n412) );
endmodule

