

module warp_checker_SHMEM_ADDR_SIZE14_DW01_cmp6_0 ( A, B, TC, LT, GT, EQ, LE, 
        GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  INV_X1 U1 ( .A(A[0]), .ZN(n3) );
  INV_X1 U2 ( .A(A[1]), .ZN(n2) );
  INV_X1 U3 ( .A(B[1]), .ZN(n1) );
  NOR4_X1 U4 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(EQ) );
  NAND4_X1 U5 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .ZN(n7) );
  XNOR2_X1 U6 ( .A(B[3]), .B(A[3]), .ZN(n11) );
  XNOR2_X1 U7 ( .A(B[4]), .B(A[4]), .ZN(n10) );
  XNOR2_X1 U8 ( .A(B[5]), .B(A[5]), .ZN(n9) );
  XNOR2_X1 U9 ( .A(B[6]), .B(A[6]), .ZN(n8) );
  NAND4_X1 U10 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .ZN(n6) );
  OAI22_X1 U11 ( .A1(n16), .A2(n2), .B1(B[1]), .B2(n16), .ZN(n15) );
  AND2_X1 U12 ( .A1(B[0]), .A2(n3), .ZN(n16) );
  OAI22_X1 U13 ( .A1(A[1]), .A2(n17), .B1(n17), .B2(n1), .ZN(n14) );
  NOR2_X1 U14 ( .A1(n3), .A2(B[0]), .ZN(n17) );
  XNOR2_X1 U15 ( .A(B[31]), .B(A[31]), .ZN(n13) );
  XNOR2_X1 U16 ( .A(B[2]), .B(A[2]), .ZN(n12) );
  NAND2_X1 U17 ( .A1(n18), .A2(n19), .ZN(n5) );
  NOR4_X1 U18 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n19) );
  XOR2_X1 U19 ( .A(B[10]), .B(A[10]), .Z(n23) );
  XOR2_X1 U20 ( .A(B[9]), .B(A[9]), .Z(n22) );
  XOR2_X1 U21 ( .A(B[8]), .B(A[8]), .Z(n21) );
  XOR2_X1 U22 ( .A(B[7]), .B(A[7]), .Z(n20) );
  NOR4_X1 U23 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n18) );
  XOR2_X1 U24 ( .A(B[14]), .B(A[14]), .Z(n27) );
  XOR2_X1 U25 ( .A(B[13]), .B(A[13]), .Z(n26) );
  XOR2_X1 U26 ( .A(B[12]), .B(A[12]), .Z(n25) );
  XOR2_X1 U27 ( .A(B[11]), .B(A[11]), .Z(n24) );
  NAND4_X1 U28 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n4) );
  NOR4_X1 U29 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(n31) );
  XOR2_X1 U30 ( .A(B[18]), .B(A[18]), .Z(n35) );
  XOR2_X1 U31 ( .A(B[17]), .B(A[17]), .Z(n34) );
  XOR2_X1 U32 ( .A(B[16]), .B(A[16]), .Z(n33) );
  XOR2_X1 U33 ( .A(B[15]), .B(A[15]), .Z(n32) );
  NOR4_X1 U34 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n30) );
  XOR2_X1 U35 ( .A(B[22]), .B(A[22]), .Z(n39) );
  XOR2_X1 U36 ( .A(B[21]), .B(A[21]), .Z(n38) );
  XOR2_X1 U37 ( .A(B[20]), .B(A[20]), .Z(n37) );
  XOR2_X1 U38 ( .A(B[19]), .B(A[19]), .Z(n36) );
  NOR4_X1 U39 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n29) );
  XOR2_X1 U40 ( .A(B[26]), .B(A[26]), .Z(n43) );
  XOR2_X1 U41 ( .A(B[25]), .B(A[25]), .Z(n42) );
  XOR2_X1 U42 ( .A(B[24]), .B(A[24]), .Z(n41) );
  XOR2_X1 U43 ( .A(B[23]), .B(A[23]), .Z(n40) );
  NOR4_X1 U44 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n28) );
  XOR2_X1 U45 ( .A(B[30]), .B(A[30]), .Z(n47) );
  XOR2_X1 U46 ( .A(B[29]), .B(A[29]), .Z(n46) );
  XOR2_X1 U47 ( .A(B[28]), .B(A[28]), .Z(n45) );
  XOR2_X1 U48 ( .A(B[27]), .B(A[27]), .Z(n44) );
endmodule


module warp_checker ( clk_in, host_reset, reset, en, 
        warp_id_in, warp_lane_id_in, cta_id_in, initial_mask_in, 
        current_mask_in, shmem_base_addr_in, gprs_base_addr_in, next_pc_in, 
        warp_state_in, warps_per_block_in, warp_pool_addr_out, 
        warp_pool_wr_en_out, warp_pool_wr_data_out, warp_state_addr_out, 
        warp_state_wr_en_out, warp_state_wr_data_out, fence_regs_fence_en_out, 
        fence_regs_fence_en_ld, .fence_regs_cta_id_in({
        \fence_regs_cta_id_in[31><3] , \fence_regs_cta_id_in[31><2] , 
        \fence_regs_cta_id_in[31><1] , \fence_regs_cta_id_in[31><0] , 
        \fence_regs_cta_id_in[30><3] , \fence_regs_cta_id_in[30><2] , 
        \fence_regs_cta_id_in[30><1] , \fence_regs_cta_id_in[30><0] , 
        \fence_regs_cta_id_in[29><3] , \fence_regs_cta_id_in[29><2] , 
        \fence_regs_cta_id_in[29><1] , \fence_regs_cta_id_in[29><0] , 
        \fence_regs_cta_id_in[28><3] , \fence_regs_cta_id_in[28><2] , 
        \fence_regs_cta_id_in[28><1] , \fence_regs_cta_id_in[28><0] , 
        \fence_regs_cta_id_in[27><3] , \fence_regs_cta_id_in[27><2] , 
        \fence_regs_cta_id_in[27><1] , \fence_regs_cta_id_in[27><0] , 
        \fence_regs_cta_id_in[26><3] , \fence_regs_cta_id_in[26><2] , 
        \fence_regs_cta_id_in[26><1] , \fence_regs_cta_id_in[26><0] , 
        \fence_regs_cta_id_in[25><3] , \fence_regs_cta_id_in[25><2] , 
        \fence_regs_cta_id_in[25><1] , \fence_regs_cta_id_in[25><0] , 
        \fence_regs_cta_id_in[24><3] , \fence_regs_cta_id_in[24><2] , 
        \fence_regs_cta_id_in[24><1] , \fence_regs_cta_id_in[24><0] , 
        \fence_regs_cta_id_in[23><3] , \fence_regs_cta_id_in[23><2] , 
        \fence_regs_cta_id_in[23><1] , \fence_regs_cta_id_in[23><0] , 
        \fence_regs_cta_id_in[22><3] , \fence_regs_cta_id_in[22><2] , 
        \fence_regs_cta_id_in[22><1] , \fence_regs_cta_id_in[22><0] , 
        \fence_regs_cta_id_in[21><3] , \fence_regs_cta_id_in[21><2] , 
        \fence_regs_cta_id_in[21><1] , \fence_regs_cta_id_in[21><0] , 
        \fence_regs_cta_id_in[20><3] , \fence_regs_cta_id_in[20><2] , 
        \fence_regs_cta_id_in[20><1] , \fence_regs_cta_id_in[20><0] , 
        \fence_regs_cta_id_in[19><3] , \fence_regs_cta_id_in[19><2] , 
        \fence_regs_cta_id_in[19><1] , \fence_regs_cta_id_in[19><0] , 
        \fence_regs_cta_id_in[18><3] , \fence_regs_cta_id_in[18><2] , 
        \fence_regs_cta_id_in[18><1] , \fence_regs_cta_id_in[18><0] , 
        \fence_regs_cta_id_in[17><3] , \fence_regs_cta_id_in[17><2] , 
        \fence_regs_cta_id_in[17><1] , \fence_regs_cta_id_in[17><0] , 
        \fence_regs_cta_id_in[16><3] , \fence_regs_cta_id_in[16><2] , 
        \fence_regs_cta_id_in[16><1] , \fence_regs_cta_id_in[16><0] , 
        \fence_regs_cta_id_in[15><3] , \fence_regs_cta_id_in[15><2] , 
        \fence_regs_cta_id_in[15><1] , \fence_regs_cta_id_in[15><0] , 
        \fence_regs_cta_id_in[14><3] , \fence_regs_cta_id_in[14><2] , 
        \fence_regs_cta_id_in[14><1] , \fence_regs_cta_id_in[14><0] , 
        \fence_regs_cta_id_in[13><3] , \fence_regs_cta_id_in[13><2] , 
        \fence_regs_cta_id_in[13><1] , \fence_regs_cta_id_in[13><0] , 
        \fence_regs_cta_id_in[12><3] , \fence_regs_cta_id_in[12><2] , 
        \fence_regs_cta_id_in[12><1] , \fence_regs_cta_id_in[12><0] , 
        \fence_regs_cta_id_in[11><3] , \fence_regs_cta_id_in[11><2] , 
        \fence_regs_cta_id_in[11><1] , \fence_regs_cta_id_in[11><0] , 
        \fence_regs_cta_id_in[10><3] , \fence_regs_cta_id_in[10><2] , 
        \fence_regs_cta_id_in[10><1] , \fence_regs_cta_id_in[10><0] , 
        \fence_regs_cta_id_in[9><3] , \fence_regs_cta_id_in[9><2] , 
        \fence_regs_cta_id_in[9><1] , \fence_regs_cta_id_in[9><0] , 
        \fence_regs_cta_id_in[8><3] , \fence_regs_cta_id_in[8><2] , 
        \fence_regs_cta_id_in[8><1] , \fence_regs_cta_id_in[8><0] , 
        \fence_regs_cta_id_in[7><3] , \fence_regs_cta_id_in[7><2] , 
        \fence_regs_cta_id_in[7><1] , \fence_regs_cta_id_in[7><0] , 
        \fence_regs_cta_id_in[6><3] , \fence_regs_cta_id_in[6><2] , 
        \fence_regs_cta_id_in[6><1] , \fence_regs_cta_id_in[6><0] , 
        \fence_regs_cta_id_in[5><3] , \fence_regs_cta_id_in[5><2] , 
        \fence_regs_cta_id_in[5><1] , \fence_regs_cta_id_in[5><0] , 
        \fence_regs_cta_id_in[4><3] , \fence_regs_cta_id_in[4><2] , 
        \fence_regs_cta_id_in[4><1] , \fence_regs_cta_id_in[4><0] , 
        \fence_regs_cta_id_in[3><3] , \fence_regs_cta_id_in[3><2] , 
        \fence_regs_cta_id_in[3><1] , \fence_regs_cta_id_in[3><0] , 
        \fence_regs_cta_id_in[2><3] , \fence_regs_cta_id_in[2><2] , 
        \fence_regs_cta_id_in[2><1] , \fence_regs_cta_id_in[2><0] , 
        \fence_regs_cta_id_in[1><3] , \fence_regs_cta_id_in[1><2] , 
        \fence_regs_cta_id_in[1><1] , \fence_regs_cta_id_in[1><0] , 
        \fence_regs_cta_id_in[0><3] , \fence_regs_cta_id_in[0><2] , 
        \fence_regs_cta_id_in[0><1] , \fence_regs_cta_id_in[0><0] }), 
        fence_regs_fence_en_in, warps_done_mask_out, pipeline_stall_out );
  input [4:0] warp_id_in;
  input [1:0] warp_lane_id_in;
  input [3:0] cta_id_in;
  input [31:0] initial_mask_in;
  input [31:0] current_mask_in;
  input [13:0] shmem_base_addr_in;
  input [8:0] gprs_base_addr_in;
  input [31:0] next_pc_in;
  input [1:0] warp_state_in;
  input [5:0] warps_per_block_in;
  output [4:0] warp_pool_addr_out;
  output [127:0] warp_pool_wr_data_out;
  output [4:0] warp_state_addr_out;
  output [1:0] warp_state_wr_data_out;
  output [31:0] fence_regs_fence_en_out;
  output [31:0] fence_regs_fence_en_ld;
  input [31:0] fence_regs_fence_en_in;
  output [31:0] warps_done_mask_out;
  input clk_in, host_reset, reset, en, \fence_regs_cta_id_in[31><3] ,
         \fence_regs_cta_id_in[31><2] , \fence_regs_cta_id_in[31><1] ,
         \fence_regs_cta_id_in[31><0] , \fence_regs_cta_id_in[30><3] ,
         \fence_regs_cta_id_in[30><2] , \fence_regs_cta_id_in[30><1] ,
         \fence_regs_cta_id_in[30><0] , \fence_regs_cta_id_in[29><3] ,
         \fence_regs_cta_id_in[29><2] , \fence_regs_cta_id_in[29><1] ,
         \fence_regs_cta_id_in[29><0] , \fence_regs_cta_id_in[28><3] ,
         \fence_regs_cta_id_in[28><2] , \fence_regs_cta_id_in[28><1] ,
         \fence_regs_cta_id_in[28><0] , \fence_regs_cta_id_in[27><3] ,
         \fence_regs_cta_id_in[27><2] , \fence_regs_cta_id_in[27><1] ,
         \fence_regs_cta_id_in[27><0] , \fence_regs_cta_id_in[26><3] ,
         \fence_regs_cta_id_in[26><2] , \fence_regs_cta_id_in[26><1] ,
         \fence_regs_cta_id_in[26><0] , \fence_regs_cta_id_in[25><3] ,
         \fence_regs_cta_id_in[25><2] , \fence_regs_cta_id_in[25><1] ,
         \fence_regs_cta_id_in[25><0] , \fence_regs_cta_id_in[24><3] ,
         \fence_regs_cta_id_in[24><2] , \fence_regs_cta_id_in[24><1] ,
         \fence_regs_cta_id_in[24><0] , \fence_regs_cta_id_in[23><3] ,
         \fence_regs_cta_id_in[23><2] , \fence_regs_cta_id_in[23><1] ,
         \fence_regs_cta_id_in[23><0] , \fence_regs_cta_id_in[22><3] ,
         \fence_regs_cta_id_in[22><2] , \fence_regs_cta_id_in[22><1] ,
         \fence_regs_cta_id_in[22><0] , \fence_regs_cta_id_in[21><3] ,
         \fence_regs_cta_id_in[21><2] , \fence_regs_cta_id_in[21><1] ,
         \fence_regs_cta_id_in[21><0] , \fence_regs_cta_id_in[20><3] ,
         \fence_regs_cta_id_in[20><2] , \fence_regs_cta_id_in[20><1] ,
         \fence_regs_cta_id_in[20><0] , \fence_regs_cta_id_in[19><3] ,
         \fence_regs_cta_id_in[19><2] , \fence_regs_cta_id_in[19><1] ,
         \fence_regs_cta_id_in[19><0] , \fence_regs_cta_id_in[18><3] ,
         \fence_regs_cta_id_in[18><2] , \fence_regs_cta_id_in[18><1] ,
         \fence_regs_cta_id_in[18><0] , \fence_regs_cta_id_in[17><3] ,
         \fence_regs_cta_id_in[17><2] , \fence_regs_cta_id_in[17><1] ,
         \fence_regs_cta_id_in[17><0] , \fence_regs_cta_id_in[16><3] ,
         \fence_regs_cta_id_in[16><2] , \fence_regs_cta_id_in[16><1] ,
         \fence_regs_cta_id_in[16><0] , \fence_regs_cta_id_in[15><3] ,
         \fence_regs_cta_id_in[15><2] , \fence_regs_cta_id_in[15><1] ,
         \fence_regs_cta_id_in[15><0] , \fence_regs_cta_id_in[14><3] ,
         \fence_regs_cta_id_in[14><2] , \fence_regs_cta_id_in[14><1] ,
         \fence_regs_cta_id_in[14><0] , \fence_regs_cta_id_in[13><3] ,
         \fence_regs_cta_id_in[13><2] , \fence_regs_cta_id_in[13><1] ,
         \fence_regs_cta_id_in[13><0] , \fence_regs_cta_id_in[12><3] ,
         \fence_regs_cta_id_in[12><2] , \fence_regs_cta_id_in[12><1] ,
         \fence_regs_cta_id_in[12><0] , \fence_regs_cta_id_in[11><3] ,
         \fence_regs_cta_id_in[11><2] , \fence_regs_cta_id_in[11><1] ,
         \fence_regs_cta_id_in[11><0] , \fence_regs_cta_id_in[10><3] ,
         \fence_regs_cta_id_in[10><2] , \fence_regs_cta_id_in[10><1] ,
         \fence_regs_cta_id_in[10><0] , \fence_regs_cta_id_in[9><3] ,
         \fence_regs_cta_id_in[9><2] , \fence_regs_cta_id_in[9><1] ,
         \fence_regs_cta_id_in[9><0] , \fence_regs_cta_id_in[8><3] ,
         \fence_regs_cta_id_in[8><2] , \fence_regs_cta_id_in[8><1] ,
         \fence_regs_cta_id_in[8><0] , \fence_regs_cta_id_in[7><3] ,
         \fence_regs_cta_id_in[7><2] , \fence_regs_cta_id_in[7><1] ,
         \fence_regs_cta_id_in[7><0] , \fence_regs_cta_id_in[6><3] ,
         \fence_regs_cta_id_in[6><2] , \fence_regs_cta_id_in[6><1] ,
         \fence_regs_cta_id_in[6><0] , \fence_regs_cta_id_in[5><3] ,
         \fence_regs_cta_id_in[5><2] , \fence_regs_cta_id_in[5><1] ,
         \fence_regs_cta_id_in[5><0] , \fence_regs_cta_id_in[4><3] ,
         \fence_regs_cta_id_in[4><2] , \fence_regs_cta_id_in[4><1] ,
         \fence_regs_cta_id_in[4><0] , \fence_regs_cta_id_in[3><3] ,
         \fence_regs_cta_id_in[3><2] , \fence_regs_cta_id_in[3><1] ,
         \fence_regs_cta_id_in[3><0] , \fence_regs_cta_id_in[2><3] ,
         \fence_regs_cta_id_in[2><2] , \fence_regs_cta_id_in[2><1] ,
         \fence_regs_cta_id_in[2><0] , \fence_regs_cta_id_in[1><3] ,
         \fence_regs_cta_id_in[1><2] , \fence_regs_cta_id_in[1><1] ,
         \fence_regs_cta_id_in[1><0] , \fence_regs_cta_id_in[0><3] ,
         \fence_regs_cta_id_in[0><2] , \fence_regs_cta_id_in[0><1] ,
         \fence_regs_cta_id_in[0><0] ;
  output warp_pool_wr_en_out, warp_state_wr_en_out, pipeline_stall_out;
  wire   N112, N113, N114, N115, N116, \warp_cntr[5] , N567, N572, N703, N704,
         N705, N706, N707, N1190, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         \add_154/carry[5] , \add_154/carry[4] , \add_154/carry[3] ,
         \add_154/carry[2] , n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651;
  wire   [4:0] warp_id_addr;
  wire   [31:0] warps_done_mask;
  wire   [2:0] warp_checker_state_machine;
  wire   [31:0] cta_id_mask_rev;
  wire   [31:0] fence_id_mask;
  assign warp_pool_wr_data_out[127] = 1'b0;
  assign warp_pool_wr_data_out[126] = 1'b0;
  assign warp_pool_wr_data_out[125] = 1'b0;
  assign warp_pool_wr_data_out[124] = 1'b0;
  assign warp_pool_wr_data_out[96] = 1'b0;
  assign N1190 = warps_per_block_in[5];

  DFFR_X1 \warp_checker_state_machine_reg[0]  ( .D(n651), .CK(clk_in), .RN(
        n132), .Q(warp_checker_state_machine[0]), .QN(n3) );
  DFFR_X1 \warp_checker_state_machine_reg[2]  ( .D(n1267), .CK(clk_in), .RN(
        n132), .Q(warp_checker_state_machine[2]), .QN(n8) );
  DFFR_X1 \warp_cntr_reg[5]  ( .D(n983), .CK(clk_in), .RN(n132), .Q(
        \warp_cntr[5] ), .QN(n9) );
  DFFR_X1 \warp_cntr_reg[4]  ( .D(n1261), .CK(clk_in), .RN(n132), .Q(N116), 
        .QN(n985) );
  DFFR_X1 \warp_checker_state_machine_reg[1]  ( .D(n1266), .CK(clk_in), .RN(
        n131), .Q(warp_checker_state_machine[1]), .QN(n7) );
  DFFR_X1 \warp_cntr_reg[3]  ( .D(n1262), .CK(clk_in), .RN(n131), .Q(N115), 
        .QN(n986) );
  DFFR_X1 \warp_cntr_reg[2]  ( .D(n1263), .CK(clk_in), .RN(n131), .Q(N114), 
        .QN(n987) );
  DFFR_X1 \warp_cntr_reg[0]  ( .D(n1264), .CK(clk_in), .RN(n131), .Q(N112), 
        .QN(n989) );
  DFFR_X1 \warp_cntr_reg[1]  ( .D(n1265), .CK(clk_in), .RN(n131), .Q(N113), 
        .QN(n988) );
  DFFR_X1 \warps_done_mask_reg[31]  ( .D(n981), .CK(clk_in), .RN(n131), .Q(
        warps_done_mask[31]), .QN(n10) );
  DFFR_X1 \warps_done_mask_reg[30]  ( .D(n980), .CK(clk_in), .RN(n131), .Q(
        warps_done_mask[30]), .QN(n11) );
  DFFR_X1 \warps_done_mask_reg[29]  ( .D(n979), .CK(clk_in), .RN(n131), .Q(
        warps_done_mask[29]), .QN(n12) );
  DFFR_X1 \warps_done_mask_reg[28]  ( .D(n978), .CK(clk_in), .RN(n131), .Q(
        warps_done_mask[28]), .QN(n13) );
  DFFR_X1 \warps_done_mask_reg[27]  ( .D(n977), .CK(clk_in), .RN(n131), .Q(
        warps_done_mask[27]), .QN(n14) );
  DFFR_X1 \warps_done_mask_reg[26]  ( .D(n976), .CK(clk_in), .RN(n131), .Q(
        warps_done_mask[26]), .QN(n15) );
  DFFR_X1 \warps_done_mask_reg[25]  ( .D(n975), .CK(clk_in), .RN(n131), .Q(
        warps_done_mask[25]), .QN(n16) );
  DFFR_X1 \warps_done_mask_reg[24]  ( .D(n974), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[24]), .QN(n17) );
  DFFR_X1 \warps_done_mask_reg[23]  ( .D(n973), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[23]), .QN(n18) );
  DFFR_X1 \warps_done_mask_reg[22]  ( .D(n972), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[22]), .QN(n19) );
  DFFR_X1 \warps_done_mask_reg[21]  ( .D(n971), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[21]), .QN(n20) );
  DFFR_X1 \warps_done_mask_reg[20]  ( .D(n970), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[20]), .QN(n21) );
  DFFR_X1 \warps_done_mask_reg[19]  ( .D(n969), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[19]), .QN(n22) );
  DFFR_X1 \warps_done_mask_reg[18]  ( .D(n968), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[18]), .QN(n23) );
  DFFR_X1 \warps_done_mask_reg[17]  ( .D(n967), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[17]), .QN(n24) );
  DFFR_X1 \warps_done_mask_reg[16]  ( .D(n966), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[16]), .QN(n25) );
  DFFR_X1 \warps_done_mask_reg[15]  ( .D(n965), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[15]), .QN(n26) );
  DFFR_X1 \warps_done_mask_reg[14]  ( .D(n964), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[14]), .QN(n27) );
  DFFR_X1 \warps_done_mask_reg[13]  ( .D(n963), .CK(clk_in), .RN(n130), .Q(
        warps_done_mask[13]), .QN(n28) );
  DFFR_X1 \warps_done_mask_reg[12]  ( .D(n962), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[12]), .QN(n29) );
  DFFR_X1 \warps_done_mask_reg[11]  ( .D(n961), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[11]), .QN(n30) );
  DFFR_X1 \warps_done_mask_reg[10]  ( .D(n960), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[10]), .QN(n31) );
  DFFR_X1 \warps_done_mask_reg[9]  ( .D(n959), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[9]), .QN(n32) );
  DFFR_X1 \warps_done_mask_reg[8]  ( .D(n958), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[8]), .QN(n33) );
  DFFR_X1 \warps_done_mask_reg[7]  ( .D(n957), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[7]), .QN(n34) );
  DFFR_X1 \warps_done_mask_reg[6]  ( .D(n956), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[6]), .QN(n35) );
  DFFR_X1 \warps_done_mask_reg[5]  ( .D(n955), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[5]), .QN(n36) );
  DFFR_X1 \warps_done_mask_reg[4]  ( .D(n954), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[4]), .QN(n37) );
  DFFR_X1 \warps_done_mask_reg[3]  ( .D(n953), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[3]), .QN(n38) );
  DFFR_X1 \warps_done_mask_reg[2]  ( .D(n952), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[2]), .QN(n39) );
  DFFR_X1 \warps_done_mask_reg[1]  ( .D(n951), .CK(clk_in), .RN(n129), .Q(
        warps_done_mask[1]), .QN(n40) );
  DFFR_X1 \warps_done_mask_reg[0]  ( .D(n950), .CK(clk_in), .RN(n128), .Q(
        warps_done_mask[0]), .QN(n41) );
  DFFR_X1 \fence_regs_fence_en_out_reg[16]  ( .D(n1189), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[16]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[17]  ( .D(n1190), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[17]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[18]  ( .D(n1191), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[18]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[19]  ( .D(n1192), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[19]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[20]  ( .D(n1193), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[20]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[21]  ( .D(n1194), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[21]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[22]  ( .D(n1195), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[22]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[23]  ( .D(n1196), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[23]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[24]  ( .D(n1197), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[24]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[25]  ( .D(n1198), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[25]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[26]  ( .D(n1199), .CK(clk_in), .RN(n128), .Q(fence_regs_fence_en_out[26]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[27]  ( .D(n1200), .CK(clk_in), .RN(n127), .Q(fence_regs_fence_en_out[27]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[28]  ( .D(n1201), .CK(clk_in), .RN(n127), .Q(fence_regs_fence_en_out[28]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[29]  ( .D(n1202), .CK(clk_in), .RN(n127), .Q(fence_regs_fence_en_out[29]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[30]  ( .D(n1203), .CK(clk_in), .RN(n127), .Q(fence_regs_fence_en_out[30]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[31]  ( .D(n1204), .CK(clk_in), .RN(n127), .Q(fence_regs_fence_en_out[31]) );
  DFFR_X1 \warp_id_addr_reg[1]  ( .D(n1256), .CK(clk_in), .RN(n127), .Q(
        warp_id_addr[1]), .QN(n5) );
  DFFR_X1 \warp_id_addr_reg[2]  ( .D(n1257), .CK(clk_in), .RN(n127), .Q(
        warp_id_addr[2]) );
  DFFR_X1 \warp_id_addr_reg[3]  ( .D(n1258), .CK(clk_in), .RN(n127), .Q(
        warp_id_addr[3]), .QN(n6) );
  DFFR_X1 \warp_id_addr_reg[4]  ( .D(n1259), .CK(clk_in), .RN(n127), .Q(
        warp_id_addr[4]) );
  DFFR_X1 \warp_id_addr_reg[0]  ( .D(n1260), .CK(clk_in), .RN(n127), .Q(
        warp_id_addr[0]), .QN(n4) );
  DFFR_X1 pipeline_stall_out_reg ( .D(n1255), .CK(clk_in), .RN(n127), .Q(
        pipeline_stall_out) );
  DFFR_X1 \warps_done_mask_out_reg[31]  ( .D(n1109), .CK(clk_in), .RN(n127), 
        .Q(warps_done_mask_out[31]) );
  DFFR_X1 \warps_done_mask_out_reg[30]  ( .D(n1110), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[30]) );
  DFFR_X1 \warps_done_mask_out_reg[29]  ( .D(n1111), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[29]) );
  DFFR_X1 \warps_done_mask_out_reg[28]  ( .D(n1112), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[28]) );
  DFFR_X1 \warps_done_mask_out_reg[27]  ( .D(n1113), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[27]) );
  DFFR_X1 \warps_done_mask_out_reg[26]  ( .D(n1114), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[26]) );
  DFFR_X1 \warps_done_mask_out_reg[25]  ( .D(n1115), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[25]) );
  DFFR_X1 \warps_done_mask_out_reg[24]  ( .D(n1116), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[24]) );
  DFFR_X1 \warps_done_mask_out_reg[23]  ( .D(n1117), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[23]) );
  DFFR_X1 \warps_done_mask_out_reg[22]  ( .D(n1118), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[22]) );
  DFFR_X1 \warps_done_mask_out_reg[21]  ( .D(n1119), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[21]) );
  DFFR_X1 \warps_done_mask_out_reg[20]  ( .D(n1120), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[20]) );
  DFFR_X1 \warps_done_mask_out_reg[19]  ( .D(n1121), .CK(clk_in), .RN(n126), 
        .Q(warps_done_mask_out[19]) );
  DFFR_X1 \warps_done_mask_out_reg[18]  ( .D(n1122), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[18]) );
  DFFR_X1 \warps_done_mask_out_reg[17]  ( .D(n1123), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[17]) );
  DFFR_X1 \warps_done_mask_out_reg[16]  ( .D(n1124), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[16]) );
  DFFR_X1 \warps_done_mask_out_reg[15]  ( .D(n1125), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[15]) );
  DFFR_X1 \warps_done_mask_out_reg[14]  ( .D(n1126), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[14]) );
  DFFR_X1 \warps_done_mask_out_reg[13]  ( .D(n1127), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[13]) );
  DFFR_X1 \warps_done_mask_out_reg[12]  ( .D(n1128), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[12]) );
  DFFR_X1 \warps_done_mask_out_reg[11]  ( .D(n1129), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[11]) );
  DFFR_X1 \warps_done_mask_out_reg[10]  ( .D(n1130), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[10]) );
  DFFR_X1 \warps_done_mask_out_reg[9]  ( .D(n1131), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[9]) );
  DFFR_X1 \warps_done_mask_out_reg[8]  ( .D(n1132), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[8]) );
  DFFR_X1 \warps_done_mask_out_reg[7]  ( .D(n1133), .CK(clk_in), .RN(n125), 
        .Q(warps_done_mask_out[7]) );
  DFFR_X1 \warps_done_mask_out_reg[6]  ( .D(n1134), .CK(clk_in), .RN(n124), 
        .Q(warps_done_mask_out[6]) );
  DFFR_X1 \warps_done_mask_out_reg[5]  ( .D(n1135), .CK(clk_in), .RN(n124), 
        .Q(warps_done_mask_out[5]) );
  DFFR_X1 \warps_done_mask_out_reg[4]  ( .D(n1136), .CK(clk_in), .RN(n124), 
        .Q(warps_done_mask_out[4]) );
  DFFR_X1 \warps_done_mask_out_reg[3]  ( .D(n1137), .CK(clk_in), .RN(n124), 
        .Q(warps_done_mask_out[3]) );
  DFFR_X1 \warps_done_mask_out_reg[2]  ( .D(n1138), .CK(clk_in), .RN(n124), 
        .Q(warps_done_mask_out[2]) );
  DFFR_X1 \warps_done_mask_out_reg[1]  ( .D(n1139), .CK(clk_in), .RN(n124), 
        .Q(warps_done_mask_out[1]) );
  DFFR_X1 \warps_done_mask_out_reg[0]  ( .D(n1140), .CK(clk_in), .RN(n124), 
        .Q(warps_done_mask_out[0]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[23]  ( .D(n1231), .CK(clk_in), .RN(n124), 
        .Q(fence_regs_fence_en_ld[23]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[22]  ( .D(n1232), .CK(clk_in), .RN(n124), 
        .Q(fence_regs_fence_en_ld[22]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[21]  ( .D(n1233), .CK(clk_in), .RN(n124), 
        .Q(fence_regs_fence_en_ld[21]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[20]  ( .D(n1234), .CK(clk_in), .RN(n124), 
        .Q(fence_regs_fence_en_ld[20]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[19]  ( .D(n1235), .CK(clk_in), .RN(n124), 
        .Q(fence_regs_fence_en_ld[19]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[18]  ( .D(n1236), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[18]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[17]  ( .D(n1237), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[17]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[16]  ( .D(n1238), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[16]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[31]  ( .D(n1223), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[31]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[30]  ( .D(n1224), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[30]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[29]  ( .D(n1225), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[29]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[28]  ( .D(n1226), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[28]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[27]  ( .D(n1227), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[27]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[26]  ( .D(n1228), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[26]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[25]  ( .D(n1229), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[25]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[24]  ( .D(n1230), .CK(clk_in), .RN(n123), 
        .Q(fence_regs_fence_en_ld[24]) );
  DFFR_X1 warp_pool_wr_en_out_reg ( .D(n1216), .CK(clk_in), .RN(n123), .Q(
        warp_pool_wr_en_out), .QN(n787) );
  DFFR_X1 \warp_pool_addr_out_reg[2]  ( .D(n1213), .CK(clk_in), .RN(n122), .Q(
        warp_pool_addr_out[2]), .QN(n790) );
  DFFR_X1 \warp_pool_addr_out_reg[3]  ( .D(n1214), .CK(clk_in), .RN(n122), .Q(
        warp_pool_addr_out[3]), .QN(n789) );
  DFFR_X1 \warp_pool_addr_out_reg[4]  ( .D(n1215), .CK(clk_in), .RN(n122), .Q(
        warp_pool_addr_out[4]), .QN(n788) );
  DFFR_X1 \warp_pool_addr_out_reg[1]  ( .D(n1217), .CK(clk_in), .RN(n122), .Q(
        warp_pool_addr_out[1]), .QN(n786) );
  DFFR_X1 \warp_pool_wr_data_out_reg[106]  ( .D(n1218), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[106]), .QN(n785) );
  DFFR_X1 \warp_pool_wr_data_out_reg[107]  ( .D(n1219), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[107]), .QN(n784) );
  DFFR_X1 \warp_pool_wr_data_out_reg[108]  ( .D(n1220), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[108]), .QN(n783) );
  DFFR_X1 \warp_pool_wr_data_out_reg[109]  ( .D(n1221), .CK(clk_in), .RN(n122), 
        .Q(warp_pool_wr_data_out[109]), .QN(n782) );
  DFFR_X1 \warp_pool_addr_out_reg[0]  ( .D(n1222), .CK(clk_in), .RN(n122), .Q(
        warp_pool_addr_out[0]), .QN(n781) );
  DFFR_X1 warp_state_wr_en_out_reg ( .D(n1206), .CK(clk_in), .RN(n122), .Q(
        warp_state_wr_en_out), .QN(n796) );
  DFFR_X1 \warp_state_addr_out_reg[1]  ( .D(n1207), .CK(clk_in), .RN(n122), 
        .Q(warp_state_addr_out[1]), .QN(n795) );
  DFFR_X1 \warp_state_addr_out_reg[2]  ( .D(n1208), .CK(clk_in), .RN(n122), 
        .Q(warp_state_addr_out[2]), .QN(n794) );
  DFFR_X1 \warp_state_addr_out_reg[3]  ( .D(n1209), .CK(clk_in), .RN(n121), 
        .Q(warp_state_addr_out[3]), .QN(n793) );
  DFFR_X1 \warp_state_wr_data_out_reg[0]  ( .D(n1211), .CK(clk_in), .RN(n121), 
        .Q(warp_state_wr_data_out[0]), .QN(n1173) );
  DFFR_X1 \warp_state_addr_out_reg[0]  ( .D(n1212), .CK(clk_in), .RN(n121), 
        .Q(warp_state_addr_out[0]), .QN(n791) );
  DFFR_X1 \warp_state_wr_data_out_reg[1]  ( .D(n984), .CK(clk_in), .RN(n121), 
        .Q(warp_state_wr_data_out[1]), .QN(n917) );
  DFFR_X1 \warp_pool_wr_data_out_reg[0]  ( .D(n1108), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[0]), .QN(n916) );
  DFFR_X1 \warp_pool_wr_data_out_reg[1]  ( .D(n1107), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[1]), .QN(n915) );
  DFFR_X1 \warp_pool_wr_data_out_reg[2]  ( .D(n1106), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[2]), .QN(n914) );
  DFFR_X1 \warp_pool_wr_data_out_reg[3]  ( .D(n1105), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[3]), .QN(n913) );
  DFFR_X1 \warp_pool_wr_data_out_reg[4]  ( .D(n1104), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[4]), .QN(n912) );
  DFFR_X1 \warp_pool_wr_data_out_reg[5]  ( .D(n1103), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[5]), .QN(n911) );
  DFFR_X1 \warp_pool_wr_data_out_reg[6]  ( .D(n1102), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[6]), .QN(n910) );
  DFFR_X1 \warp_pool_wr_data_out_reg[7]  ( .D(n1101), .CK(clk_in), .RN(n121), 
        .Q(warp_pool_wr_data_out[7]), .QN(n909) );
  DFFR_X1 \warp_pool_wr_data_out_reg[8]  ( .D(n1100), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[8]), .QN(n908) );
  DFFR_X1 \warp_pool_wr_data_out_reg[9]  ( .D(n1099), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[9]), .QN(n907) );
  DFFR_X1 \warp_pool_wr_data_out_reg[10]  ( .D(n1098), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[10]), .QN(n906) );
  DFFR_X1 \warp_pool_wr_data_out_reg[11]  ( .D(n1097), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[11]), .QN(n905) );
  DFFR_X1 \warp_pool_wr_data_out_reg[12]  ( .D(n1096), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[12]), .QN(n904) );
  DFFR_X1 \warp_pool_wr_data_out_reg[13]  ( .D(n1095), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[13]), .QN(n903) );
  DFFR_X1 \warp_pool_wr_data_out_reg[14]  ( .D(n1094), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[14]), .QN(n902) );
  DFFR_X1 \warp_pool_wr_data_out_reg[15]  ( .D(n1093), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[15]), .QN(n901) );
  DFFR_X1 \warp_pool_wr_data_out_reg[16]  ( .D(n1092), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[16]), .QN(n900) );
  DFFR_X1 \warp_pool_wr_data_out_reg[17]  ( .D(n1091), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[17]), .QN(n899) );
  DFFR_X1 \warp_pool_wr_data_out_reg[18]  ( .D(n1090), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[18]), .QN(n898) );
  DFFR_X1 \warp_pool_wr_data_out_reg[19]  ( .D(n1089), .CK(clk_in), .RN(n120), 
        .Q(warp_pool_wr_data_out[19]), .QN(n897) );
  DFFR_X1 \warp_pool_wr_data_out_reg[20]  ( .D(n1088), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[20]), .QN(n896) );
  DFFR_X1 \warp_pool_wr_data_out_reg[21]  ( .D(n1087), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[21]), .QN(n895) );
  DFFR_X1 \warp_pool_wr_data_out_reg[22]  ( .D(n1086), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[22]), .QN(n894) );
  DFFR_X1 \warp_pool_wr_data_out_reg[23]  ( .D(n1085), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[23]), .QN(n893) );
  DFFR_X1 \warp_pool_wr_data_out_reg[24]  ( .D(n1084), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[24]), .QN(n892) );
  DFFR_X1 \warp_pool_wr_data_out_reg[25]  ( .D(n1083), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[25]), .QN(n891) );
  DFFR_X1 \warp_pool_wr_data_out_reg[26]  ( .D(n1082), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[26]), .QN(n890) );
  DFFR_X1 \warp_pool_wr_data_out_reg[27]  ( .D(n1081), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[27]), .QN(n889) );
  DFFR_X1 \warp_pool_wr_data_out_reg[28]  ( .D(n1080), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[28]), .QN(n888) );
  DFFR_X1 \warp_pool_wr_data_out_reg[29]  ( .D(n1079), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[29]), .QN(n887) );
  DFFR_X1 \warp_pool_wr_data_out_reg[30]  ( .D(n1078), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[30]), .QN(n886) );
  DFFR_X1 \warp_pool_wr_data_out_reg[31]  ( .D(n1077), .CK(clk_in), .RN(n119), 
        .Q(warp_pool_wr_data_out[31]), .QN(n885) );
  DFFR_X1 \warp_pool_wr_data_out_reg[32]  ( .D(n1076), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[32]), .QN(n884) );
  DFFR_X1 \warp_pool_wr_data_out_reg[33]  ( .D(n1075), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[33]), .QN(n883) );
  DFFR_X1 \warp_pool_wr_data_out_reg[34]  ( .D(n1074), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[34]), .QN(n882) );
  DFFR_X1 \warp_pool_wr_data_out_reg[35]  ( .D(n1073), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[35]), .QN(n881) );
  DFFR_X1 \warp_pool_wr_data_out_reg[36]  ( .D(n1072), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[36]), .QN(n880) );
  DFFR_X1 \warp_pool_wr_data_out_reg[37]  ( .D(n1071), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[37]), .QN(n879) );
  DFFR_X1 \warp_pool_wr_data_out_reg[38]  ( .D(n1070), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[38]), .QN(n878) );
  DFFR_X1 \warp_pool_wr_data_out_reg[39]  ( .D(n1069), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[39]), .QN(n877) );
  DFFR_X1 \warp_pool_wr_data_out_reg[40]  ( .D(n1068), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[40]), .QN(n876) );
  DFFR_X1 \warp_pool_wr_data_out_reg[41]  ( .D(n1067), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[41]), .QN(n875) );
  DFFR_X1 \warp_pool_wr_data_out_reg[42]  ( .D(n1066), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[42]), .QN(n874) );
  DFFR_X1 \warp_pool_wr_data_out_reg[43]  ( .D(n1065), .CK(clk_in), .RN(n118), 
        .Q(warp_pool_wr_data_out[43]), .QN(n873) );
  DFFR_X1 \warp_pool_wr_data_out_reg[44]  ( .D(n1064), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[44]), .QN(n872) );
  DFFR_X1 \warp_pool_wr_data_out_reg[45]  ( .D(n1063), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[45]), .QN(n871) );
  DFFR_X1 \warp_pool_wr_data_out_reg[46]  ( .D(n1062), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[46]), .QN(n870) );
  DFFR_X1 \warp_pool_wr_data_out_reg[47]  ( .D(n1061), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[47]), .QN(n869) );
  DFFR_X1 \warp_pool_wr_data_out_reg[48]  ( .D(n1060), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[48]), .QN(n868) );
  DFFR_X1 \warp_pool_wr_data_out_reg[49]  ( .D(n1059), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[49]), .QN(n867) );
  DFFR_X1 \warp_pool_wr_data_out_reg[50]  ( .D(n1058), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[50]), .QN(n866) );
  DFFR_X1 \warp_pool_wr_data_out_reg[51]  ( .D(n1057), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[51]), .QN(n865) );
  DFFR_X1 \warp_pool_wr_data_out_reg[52]  ( .D(n1056), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[52]), .QN(n864) );
  DFFR_X1 \warp_pool_wr_data_out_reg[53]  ( .D(n1055), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[53]), .QN(n863) );
  DFFR_X1 \warp_pool_wr_data_out_reg[54]  ( .D(n1054), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[54]), .QN(n862) );
  DFFR_X1 \warp_pool_wr_data_out_reg[55]  ( .D(n1053), .CK(clk_in), .RN(n117), 
        .Q(warp_pool_wr_data_out[55]), .QN(n861) );
  DFFR_X1 \warp_pool_wr_data_out_reg[56]  ( .D(n1052), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[56]), .QN(n860) );
  DFFR_X1 \warp_pool_wr_data_out_reg[57]  ( .D(n1051), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[57]), .QN(n859) );
  DFFR_X1 \warp_pool_wr_data_out_reg[58]  ( .D(n1050), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[58]), .QN(n858) );
  DFFR_X1 \warp_pool_wr_data_out_reg[59]  ( .D(n1049), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[59]), .QN(n857) );
  DFFR_X1 \warp_pool_wr_data_out_reg[60]  ( .D(n1048), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[60]), .QN(n856) );
  DFFR_X1 \warp_pool_wr_data_out_reg[61]  ( .D(n1047), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[61]), .QN(n855) );
  DFFR_X1 \warp_pool_wr_data_out_reg[62]  ( .D(n1046), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[62]), .QN(n854) );
  DFFR_X1 \warp_pool_wr_data_out_reg[63]  ( .D(n1045), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[63]), .QN(n853) );
  DFFR_X1 \warp_pool_wr_data_out_reg[64]  ( .D(n1044), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[64]), .QN(n852) );
  DFFR_X1 \warp_pool_wr_data_out_reg[65]  ( .D(n1043), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[65]), .QN(n851) );
  DFFR_X1 \warp_pool_wr_data_out_reg[66]  ( .D(n1042), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[66]), .QN(n850) );
  DFFR_X1 \warp_pool_wr_data_out_reg[67]  ( .D(n1041), .CK(clk_in), .RN(n116), 
        .Q(warp_pool_wr_data_out[67]), .QN(n849) );
  DFFR_X1 \warp_pool_wr_data_out_reg[68]  ( .D(n1040), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[68]), .QN(n848) );
  DFFR_X1 \warp_pool_wr_data_out_reg[69]  ( .D(n1039), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[69]), .QN(n847) );
  DFFR_X1 \warp_pool_wr_data_out_reg[70]  ( .D(n1038), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[70]), .QN(n846) );
  DFFR_X1 \warp_pool_wr_data_out_reg[71]  ( .D(n1037), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[71]), .QN(n845) );
  DFFR_X1 \warp_pool_wr_data_out_reg[72]  ( .D(n1036), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[72]), .QN(n844) );
  DFFR_X1 \warp_pool_wr_data_out_reg[73]  ( .D(n1035), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[73]), .QN(n843) );
  DFFR_X1 \warp_pool_wr_data_out_reg[74]  ( .D(n1034), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[74]), .QN(n842) );
  DFFR_X1 \warp_pool_wr_data_out_reg[75]  ( .D(n1033), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[75]), .QN(n841) );
  DFFR_X1 \warp_pool_wr_data_out_reg[76]  ( .D(n1032), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[76]), .QN(n840) );
  DFFR_X1 \warp_pool_wr_data_out_reg[77]  ( .D(n1031), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[77]), .QN(n839) );
  DFFR_X1 \warp_pool_wr_data_out_reg[78]  ( .D(n1030), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[78]), .QN(n838) );
  DFFR_X1 \warp_pool_wr_data_out_reg[79]  ( .D(n1029), .CK(clk_in), .RN(n115), 
        .Q(warp_pool_wr_data_out[79]), .QN(n837) );
  DFFR_X1 \warp_pool_wr_data_out_reg[80]  ( .D(n1028), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[80]), .QN(n836) );
  DFFR_X1 \warp_pool_wr_data_out_reg[81]  ( .D(n1027), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[81]), .QN(n835) );
  DFFR_X1 \warp_pool_wr_data_out_reg[82]  ( .D(n1026), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[82]), .QN(n834) );
  DFFR_X1 \warp_pool_wr_data_out_reg[83]  ( .D(n1025), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[83]), .QN(n833) );
  DFFR_X1 \warp_pool_wr_data_out_reg[84]  ( .D(n1024), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[84]), .QN(n832) );
  DFFR_X1 \warp_pool_wr_data_out_reg[85]  ( .D(n1023), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[85]), .QN(n831) );
  DFFR_X1 \warp_pool_wr_data_out_reg[86]  ( .D(n1022), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[86]), .QN(n830) );
  DFFR_X1 \warp_pool_wr_data_out_reg[87]  ( .D(n1021), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[87]), .QN(n829) );
  DFFR_X1 \warp_pool_wr_data_out_reg[88]  ( .D(n1020), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[88]), .QN(n828) );
  DFFR_X1 \warp_pool_wr_data_out_reg[89]  ( .D(n1019), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[89]), .QN(n827) );
  DFFR_X1 \warp_pool_wr_data_out_reg[90]  ( .D(n1018), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[90]), .QN(n826) );
  DFFR_X1 \warp_pool_wr_data_out_reg[91]  ( .D(n1017), .CK(clk_in), .RN(n114), 
        .Q(warp_pool_wr_data_out[91]), .QN(n825) );
  DFFR_X1 \warp_pool_wr_data_out_reg[92]  ( .D(n1016), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[92]), .QN(n824) );
  DFFR_X1 \warp_pool_wr_data_out_reg[93]  ( .D(n1015), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[93]), .QN(n823) );
  DFFR_X1 \warp_pool_wr_data_out_reg[94]  ( .D(n1014), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[94]), .QN(n822) );
  DFFR_X1 \warp_pool_wr_data_out_reg[95]  ( .D(n1013), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[95]), .QN(n821) );
  DFFR_X1 \warp_pool_wr_data_out_reg[97]  ( .D(n1012), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[97]), .QN(n820) );
  DFFR_X1 \warp_pool_wr_data_out_reg[98]  ( .D(n1011), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[98]), .QN(n819) );
  DFFR_X1 \warp_pool_wr_data_out_reg[99]  ( .D(n1010), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[99]), .QN(n818) );
  DFFR_X1 \warp_pool_wr_data_out_reg[100]  ( .D(n1009), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[100]), .QN(n817) );
  DFFR_X1 \warp_pool_wr_data_out_reg[101]  ( .D(n1008), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[101]), .QN(n816) );
  DFFR_X1 \warp_pool_wr_data_out_reg[102]  ( .D(n1007), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[102]), .QN(n815) );
  DFFR_X1 \warp_pool_wr_data_out_reg[103]  ( .D(n1006), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[103]), .QN(n814) );
  DFFR_X1 \warp_pool_wr_data_out_reg[104]  ( .D(n1005), .CK(clk_in), .RN(n113), 
        .Q(warp_pool_wr_data_out[104]), .QN(n813) );
  DFFR_X1 \warp_pool_wr_data_out_reg[105]  ( .D(n1004), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[105]), .QN(n812) );
  DFFR_X1 \warp_pool_wr_data_out_reg[110]  ( .D(n1003), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[110]), .QN(n811) );
  DFFR_X1 \warp_pool_wr_data_out_reg[111]  ( .D(n1002), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[111]), .QN(n810) );
  DFFR_X1 \warp_pool_wr_data_out_reg[112]  ( .D(n1001), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[112]), .QN(n809) );
  DFFR_X1 \warp_pool_wr_data_out_reg[113]  ( .D(n1000), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[113]), .QN(n808) );
  DFFR_X1 \warp_pool_wr_data_out_reg[114]  ( .D(n999), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[114]), .QN(n807) );
  DFFR_X1 \warp_pool_wr_data_out_reg[115]  ( .D(n998), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[115]), .QN(n806) );
  DFFR_X1 \warp_pool_wr_data_out_reg[116]  ( .D(n997), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[116]), .QN(n805) );
  DFFR_X1 \warp_pool_wr_data_out_reg[117]  ( .D(n996), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[117]), .QN(n804) );
  DFFR_X1 \warp_pool_wr_data_out_reg[118]  ( .D(n995), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[118]), .QN(n803) );
  DFFR_X1 \warp_pool_wr_data_out_reg[119]  ( .D(n994), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[119]), .QN(n802) );
  DFFR_X1 \warp_pool_wr_data_out_reg[120]  ( .D(n993), .CK(clk_in), .RN(n112), 
        .Q(warp_pool_wr_data_out[120]), .QN(n801) );
  DFFR_X1 \warp_pool_wr_data_out_reg[121]  ( .D(n992), .CK(clk_in), .RN(n111), 
        .Q(warp_pool_wr_data_out[121]), .QN(n800) );
  DFFR_X1 \warp_pool_wr_data_out_reg[122]  ( .D(n991), .CK(clk_in), .RN(n111), 
        .Q(warp_pool_wr_data_out[122]), .QN(n799) );
  DFFR_X1 \warp_pool_wr_data_out_reg[123]  ( .D(n990), .CK(clk_in), .RN(n111), 
        .Q(warp_pool_wr_data_out[123]), .QN(n798) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[7]  ( .D(n1247), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_ld[7]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[7]  ( .D(n1180), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_out[7]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[6]  ( .D(n1248), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_ld[6]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[6]  ( .D(n1179), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_out[6]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[5]  ( .D(n1249), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_ld[5]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[5]  ( .D(n1178), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_out[5]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[4]  ( .D(n1250), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_ld[4]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[4]  ( .D(n1177), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_out[4]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[3]  ( .D(n1251), .CK(clk_in), .RN(n111), 
        .Q(fence_regs_fence_en_ld[3]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[3]  ( .D(n1176), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_out[3]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[2]  ( .D(n1252), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_ld[2]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[2]  ( .D(n1175), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_out[2]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[1]  ( .D(n1253), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_ld[1]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[1]  ( .D(n1174), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_out[1]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[0]  ( .D(n1254), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_ld[0]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[0]  ( .D(n1205), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_out[0]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[15]  ( .D(n1239), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_ld[15]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[15]  ( .D(n1188), .CK(clk_in), .RN(n110), .Q(fence_regs_fence_en_out[15]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[14]  ( .D(n1240), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_ld[14]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[14]  ( .D(n1187), .CK(clk_in), .RN(n110), .Q(fence_regs_fence_en_out[14]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[13]  ( .D(n1241), .CK(clk_in), .RN(n110), 
        .Q(fence_regs_fence_en_ld[13]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[13]  ( .D(n1186), .CK(clk_in), .RN(n109), .Q(fence_regs_fence_en_out[13]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[12]  ( .D(n1242), .CK(clk_in), .RN(n109), 
        .Q(fence_regs_fence_en_ld[12]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[12]  ( .D(n1185), .CK(clk_in), .RN(n109), .Q(fence_regs_fence_en_out[12]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[11]  ( .D(n1243), .CK(clk_in), .RN(n109), 
        .Q(fence_regs_fence_en_ld[11]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[11]  ( .D(n1184), .CK(clk_in), .RN(n109), .Q(fence_regs_fence_en_out[11]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[10]  ( .D(n1244), .CK(clk_in), .RN(n109), 
        .Q(fence_regs_fence_en_ld[10]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[10]  ( .D(n1183), .CK(clk_in), .RN(n109), .Q(fence_regs_fence_en_out[10]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[9]  ( .D(n1245), .CK(clk_in), .RN(n109), 
        .Q(fence_regs_fence_en_ld[9]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[9]  ( .D(n1182), .CK(clk_in), .RN(n109), 
        .Q(fence_regs_fence_en_out[9]) );
  DFFR_X1 \fence_regs_fence_en_ld_reg[8]  ( .D(n1246), .CK(clk_in), .RN(n109), 
        .Q(fence_regs_fence_en_ld[8]) );
  DFFR_X1 \fence_regs_fence_en_out_reg[8]  ( .D(n1181), .CK(clk_in), .RN(n109), 
        .Q(fence_regs_fence_en_out[8]) );
  DFFR_X1 \warp_state_addr_out_reg[4]  ( .D(n1210), .CK(clk_in), .RN(n109), 
        .Q(warp_state_addr_out[4]), .QN(n792) );
  warp_checker_SHMEM_ADDR_SIZE14_DW01_cmp6_0 eq_137 ( .A(cta_id_mask_rev), .B(
        fence_id_mask), .TC(1'b0), .EQ(N567) );
  HA_X1 \add_154/U1_1_1  ( .A(N113), .B(N112), .CO(\add_154/carry[2] ), .S(
        N703) );
  HA_X1 \add_154/U1_1_2  ( .A(N114), .B(\add_154/carry[2] ), .CO(
        \add_154/carry[3] ), .S(N704) );
  HA_X1 \add_154/U1_1_3  ( .A(N115), .B(\add_154/carry[3] ), .CO(
        \add_154/carry[4] ), .S(N705) );
  HA_X1 \add_154/U1_1_4  ( .A(N116), .B(\add_154/carry[4] ), .CO(
        \add_154/carry[5] ), .S(N706) );
  AND3_X1 U3 ( .A1(n197), .A2(n187), .A3(n414), .ZN(n1) );
  NOR3_X2 U4 ( .A1(n6), .A2(warp_id_addr[4]), .A3(n187), .ZN(n224) );
  NOR3_X2 U5 ( .A1(warp_id_addr[3]), .A2(warp_id_addr[4]), .A3(n187), .ZN(n200) );
  BUF_X1 U6 ( .A(n94), .Z(n89) );
  BUF_X1 U7 ( .A(n94), .Z(n88) );
  BUF_X1 U9 ( .A(n94), .Z(n93) );
  BUF_X1 U10 ( .A(n95), .Z(n87) );
  BUF_X1 U11 ( .A(n95), .Z(n86) );
  BUF_X1 U12 ( .A(n95), .Z(n85) );
  BUF_X1 U13 ( .A(n95), .Z(n84) );
  BUF_X1 U14 ( .A(n94), .Z(n92) );
  BUF_X1 U15 ( .A(n94), .Z(n91) );
  BUF_X1 U16 ( .A(n94), .Z(n90) );
  BUF_X1 U17 ( .A(n95), .Z(n83) );
  INV_X1 U18 ( .A(n1), .ZN(n82) );
  INV_X1 U19 ( .A(n1), .ZN(n79) );
  BUF_X1 U20 ( .A(n163), .Z(n96) );
  BUF_X1 U21 ( .A(n163), .Z(n97) );
  BUF_X1 U22 ( .A(n149), .Z(n94) );
  BUF_X1 U23 ( .A(n163), .Z(n98) );
  BUF_X1 U24 ( .A(n149), .Z(n95) );
  BUF_X1 U25 ( .A(n108), .Z(n136) );
  BUF_X1 U26 ( .A(n108), .Z(n135) );
  BUF_X1 U27 ( .A(n107), .Z(n134) );
  BUF_X1 U28 ( .A(n107), .Z(n133) );
  INV_X1 U29 ( .A(n102), .ZN(n100) );
  INV_X1 U30 ( .A(n102), .ZN(n99) );
  BUF_X1 U31 ( .A(n103), .Z(n105) );
  BUF_X1 U32 ( .A(n103), .Z(n104) );
  BUF_X1 U33 ( .A(n103), .Z(n106) );
  BUF_X1 U34 ( .A(n982), .Z(n108) );
  BUF_X1 U35 ( .A(n982), .Z(n107) );
  INV_X1 U36 ( .A(n138), .ZN(n137) );
  INV_X1 U37 ( .A(n140), .ZN(n139) );
  INV_X1 U38 ( .A(n142), .ZN(n141) );
  INV_X1 U39 ( .A(n144), .ZN(n143) );
  INV_X1 U40 ( .A(n53), .ZN(n73) );
  INV_X1 U41 ( .A(n47), .ZN(n71) );
  INV_X1 U42 ( .A(n54), .ZN(n74) );
  NAND2_X1 U43 ( .A1(n1), .A2(n281), .ZN(n160) );
  INV_X1 U44 ( .A(n44), .ZN(n70) );
  INV_X1 U45 ( .A(n60), .ZN(n76) );
  INV_X1 U46 ( .A(n57), .ZN(n75) );
  BUF_X1 U47 ( .A(n42), .Z(n102) );
  BUF_X1 U48 ( .A(n42), .Z(n101) );
  BUF_X1 U49 ( .A(n303), .Z(n103) );
  INV_X1 U50 ( .A(n43), .ZN(n69) );
  INV_X1 U51 ( .A(n48), .ZN(n72) );
  INV_X1 U52 ( .A(cta_id_in[1]), .ZN(n140) );
  INV_X1 U53 ( .A(cta_id_in[3]), .ZN(n144) );
  INV_X1 U54 ( .A(cta_id_in[2]), .ZN(n142) );
  INV_X1 U55 ( .A(cta_id_in[0]), .ZN(n138) );
  OR3_X1 U56 ( .A1(warp_checker_state_machine[1]), .A2(
        warp_checker_state_machine[2]), .A3(warp_checker_state_machine[0]), 
        .ZN(n42) );
  NOR2_X1 U57 ( .A1(n988), .A2(N112), .ZN(n62) );
  NOR2_X1 U58 ( .A1(n988), .A2(n989), .ZN(n61) );
  NOR2_X1 U59 ( .A1(N112), .A2(N113), .ZN(n59) );
  NOR2_X1 U60 ( .A1(n989), .A2(N113), .ZN(n58) );
  AOI22_X1 U61 ( .A1(cta_id_mask_rev[28]), .A2(n59), .B1(cta_id_mask_rev[29]), 
        .B2(n58), .ZN(n43) );
  AOI221_X1 U62 ( .B1(cta_id_mask_rev[30]), .B2(n62), .C1(cta_id_mask_rev[31]), 
        .C2(n61), .A(n69), .ZN(n46) );
  AOI22_X1 U63 ( .A1(cta_id_mask_rev[24]), .A2(n59), .B1(cta_id_mask_rev[25]), 
        .B2(n58), .ZN(n44) );
  AOI221_X1 U64 ( .B1(cta_id_mask_rev[26]), .B2(n62), .C1(cta_id_mask_rev[27]), 
        .C2(n61), .A(n70), .ZN(n45) );
  OAI22_X1 U65 ( .A1(n987), .A2(n46), .B1(N114), .B2(n45), .ZN(n52) );
  AOI22_X1 U66 ( .A1(cta_id_mask_rev[20]), .A2(n59), .B1(cta_id_mask_rev[21]), 
        .B2(n58), .ZN(n47) );
  AOI221_X1 U67 ( .B1(cta_id_mask_rev[22]), .B2(n62), .C1(cta_id_mask_rev[23]), 
        .C2(n61), .A(n71), .ZN(n50) );
  AOI22_X1 U68 ( .A1(cta_id_mask_rev[16]), .A2(n59), .B1(cta_id_mask_rev[17]), 
        .B2(n58), .ZN(n48) );
  AOI221_X1 U69 ( .B1(cta_id_mask_rev[18]), .B2(n62), .C1(cta_id_mask_rev[19]), 
        .C2(n61), .A(n72), .ZN(n49) );
  OAI22_X1 U70 ( .A1(n50), .A2(n987), .B1(N114), .B2(n49), .ZN(n51) );
  AOI22_X1 U71 ( .A1(N115), .A2(n52), .B1(n51), .B2(n986), .ZN(n68) );
  AOI22_X1 U72 ( .A1(cta_id_mask_rev[12]), .A2(n59), .B1(cta_id_mask_rev[13]), 
        .B2(n58), .ZN(n53) );
  AOI221_X1 U73 ( .B1(cta_id_mask_rev[14]), .B2(n62), .C1(cta_id_mask_rev[15]), 
        .C2(n61), .A(n73), .ZN(n56) );
  AOI22_X1 U74 ( .A1(cta_id_mask_rev[8]), .A2(n59), .B1(cta_id_mask_rev[9]), 
        .B2(n58), .ZN(n54) );
  AOI221_X1 U75 ( .B1(cta_id_mask_rev[10]), .B2(n62), .C1(cta_id_mask_rev[11]), 
        .C2(n61), .A(n74), .ZN(n55) );
  OAI22_X1 U76 ( .A1(n987), .A2(n56), .B1(N114), .B2(n55), .ZN(n66) );
  AOI22_X1 U77 ( .A1(cta_id_mask_rev[4]), .A2(n59), .B1(cta_id_mask_rev[5]), 
        .B2(n58), .ZN(n57) );
  AOI221_X1 U78 ( .B1(cta_id_mask_rev[6]), .B2(n62), .C1(cta_id_mask_rev[7]), 
        .C2(n61), .A(n75), .ZN(n64) );
  AOI22_X1 U79 ( .A1(cta_id_mask_rev[0]), .A2(n59), .B1(cta_id_mask_rev[1]), 
        .B2(n58), .ZN(n60) );
  AOI221_X1 U80 ( .B1(cta_id_mask_rev[2]), .B2(n62), .C1(cta_id_mask_rev[3]), 
        .C2(n61), .A(n76), .ZN(n63) );
  OAI22_X1 U81 ( .A1(n987), .A2(n64), .B1(N114), .B2(n63), .ZN(n65) );
  AOI22_X1 U82 ( .A1(n66), .A2(N115), .B1(n65), .B2(n986), .ZN(n67) );
  OAI22_X1 U83 ( .A1(n68), .A2(n985), .B1(N116), .B2(n67), .ZN(N572) );
  INV_X1 U84 ( .A(n1), .ZN(n77) );
  INV_X1 U85 ( .A(n1), .ZN(n78) );
  INV_X1 U86 ( .A(n1), .ZN(n80) );
  INV_X1 U87 ( .A(n1), .ZN(n81) );
  CLKBUF_X1 U88 ( .A(n136), .Z(n109) );
  CLKBUF_X1 U89 ( .A(n136), .Z(n110) );
  CLKBUF_X1 U90 ( .A(n136), .Z(n111) );
  CLKBUF_X1 U91 ( .A(n136), .Z(n112) );
  CLKBUF_X1 U92 ( .A(n136), .Z(n113) );
  CLKBUF_X1 U93 ( .A(n136), .Z(n114) );
  CLKBUF_X1 U94 ( .A(n135), .Z(n115) );
  CLKBUF_X1 U95 ( .A(n135), .Z(n116) );
  CLKBUF_X1 U96 ( .A(n135), .Z(n117) );
  CLKBUF_X1 U97 ( .A(n135), .Z(n118) );
  CLKBUF_X1 U98 ( .A(n135), .Z(n119) );
  CLKBUF_X1 U99 ( .A(n135), .Z(n120) );
  CLKBUF_X1 U100 ( .A(n134), .Z(n121) );
  CLKBUF_X1 U101 ( .A(n134), .Z(n122) );
  CLKBUF_X1 U102 ( .A(n134), .Z(n123) );
  CLKBUF_X1 U103 ( .A(n134), .Z(n124) );
  CLKBUF_X1 U104 ( .A(n134), .Z(n125) );
  CLKBUF_X1 U105 ( .A(n134), .Z(n126) );
  CLKBUF_X1 U106 ( .A(n133), .Z(n127) );
  CLKBUF_X1 U107 ( .A(n133), .Z(n128) );
  CLKBUF_X1 U108 ( .A(n133), .Z(n129) );
  CLKBUF_X1 U109 ( .A(n133), .Z(n130) );
  CLKBUF_X1 U110 ( .A(n133), .Z(n131) );
  CLKBUF_X1 U111 ( .A(n133), .Z(n132) );
  XOR2_X1 U112 ( .A(\add_154/carry[5] ), .B(\warp_cntr[5] ), .Z(N707) );
  OAI221_X1 U113 ( .B1(n3), .B2(n145), .C1(n146), .C2(n147), .A(n148), .ZN(
        n651) );
  OAI22_X1 U114 ( .A1(n82), .A2(n807), .B1(n88), .B2(n150), .ZN(n999) );
  INV_X1 U115 ( .A(shmem_base_addr_in[4]), .ZN(n150) );
  OAI22_X1 U116 ( .A1(n79), .A2(n806), .B1(n83), .B2(n151), .ZN(n998) );
  INV_X1 U117 ( .A(shmem_base_addr_in[5]), .ZN(n151) );
  OAI22_X1 U118 ( .A1(n81), .A2(n805), .B1(n83), .B2(n152), .ZN(n997) );
  INV_X1 U119 ( .A(shmem_base_addr_in[6]), .ZN(n152) );
  OAI22_X1 U120 ( .A1(n80), .A2(n804), .B1(n83), .B2(n153), .ZN(n996) );
  INV_X1 U121 ( .A(shmem_base_addr_in[7]), .ZN(n153) );
  OAI22_X1 U122 ( .A1(n82), .A2(n803), .B1(n83), .B2(n154), .ZN(n995) );
  INV_X1 U123 ( .A(shmem_base_addr_in[8]), .ZN(n154) );
  OAI22_X1 U124 ( .A1(n82), .A2(n802), .B1(n83), .B2(n155), .ZN(n994) );
  INV_X1 U125 ( .A(shmem_base_addr_in[9]), .ZN(n155) );
  OAI22_X1 U126 ( .A1(n78), .A2(n801), .B1(n83), .B2(n156), .ZN(n993) );
  INV_X1 U127 ( .A(shmem_base_addr_in[10]), .ZN(n156) );
  OAI22_X1 U128 ( .A1(n77), .A2(n800), .B1(n83), .B2(n157), .ZN(n992) );
  INV_X1 U129 ( .A(shmem_base_addr_in[11]), .ZN(n157) );
  OAI22_X1 U130 ( .A1(n82), .A2(n799), .B1(n84), .B2(n158), .ZN(n991) );
  INV_X1 U131 ( .A(shmem_base_addr_in[12]), .ZN(n158) );
  OAI22_X1 U132 ( .A1(n79), .A2(n798), .B1(n83), .B2(n159), .ZN(n990) );
  INV_X1 U133 ( .A(shmem_base_addr_in[13]), .ZN(n159) );
  OAI22_X1 U134 ( .A1(n160), .A2(n917), .B1(n161), .B2(n162), .ZN(n984) );
  OAI21_X1 U135 ( .B1(n9), .B2(n96), .A(n164), .ZN(n983) );
  NAND2_X1 U136 ( .A1(N707), .A2(n165), .ZN(n164) );
  NOR2_X1 U137 ( .A1(reset), .A2(host_reset), .ZN(n982) );
  OAI21_X1 U138 ( .B1(n166), .B2(n167), .A(n10), .ZN(n981) );
  OAI21_X1 U139 ( .B1(n166), .B2(n168), .A(n11), .ZN(n980) );
  OAI21_X1 U140 ( .B1(n166), .B2(n169), .A(n12), .ZN(n979) );
  OAI21_X1 U141 ( .B1(n166), .B2(n170), .A(n13), .ZN(n978) );
  OAI21_X1 U142 ( .B1(n166), .B2(n171), .A(n14), .ZN(n977) );
  OAI21_X1 U143 ( .B1(n166), .B2(n172), .A(n15), .ZN(n976) );
  OAI21_X1 U144 ( .B1(n166), .B2(n173), .A(n16), .ZN(n975) );
  OAI21_X1 U145 ( .B1(n166), .B2(n174), .A(n17), .ZN(n974) );
  NAND3_X1 U146 ( .A1(warp_id_in[3]), .A2(n175), .A3(warp_id_in[4]), .ZN(n166)
         );
  OAI21_X1 U147 ( .B1(n167), .B2(n176), .A(n18), .ZN(n973) );
  OAI21_X1 U148 ( .B1(n168), .B2(n176), .A(n19), .ZN(n972) );
  OAI21_X1 U149 ( .B1(n169), .B2(n176), .A(n20), .ZN(n971) );
  OAI21_X1 U150 ( .B1(n170), .B2(n176), .A(n21), .ZN(n970) );
  OAI21_X1 U151 ( .B1(n171), .B2(n176), .A(n22), .ZN(n969) );
  OAI21_X1 U152 ( .B1(n172), .B2(n176), .A(n23), .ZN(n968) );
  OAI21_X1 U153 ( .B1(n173), .B2(n176), .A(n24), .ZN(n967) );
  OAI21_X1 U154 ( .B1(n174), .B2(n176), .A(n25), .ZN(n966) );
  NAND3_X1 U155 ( .A1(n175), .A2(n177), .A3(warp_id_in[4]), .ZN(n176) );
  OAI21_X1 U156 ( .B1(n167), .B2(n178), .A(n26), .ZN(n965) );
  OAI21_X1 U157 ( .B1(n168), .B2(n178), .A(n27), .ZN(n964) );
  OAI21_X1 U158 ( .B1(n169), .B2(n178), .A(n28), .ZN(n963) );
  OAI21_X1 U159 ( .B1(n170), .B2(n178), .A(n29), .ZN(n962) );
  OAI21_X1 U160 ( .B1(n171), .B2(n178), .A(n30), .ZN(n961) );
  OAI21_X1 U161 ( .B1(n172), .B2(n178), .A(n31), .ZN(n960) );
  OAI21_X1 U162 ( .B1(n173), .B2(n178), .A(n32), .ZN(n959) );
  OAI21_X1 U163 ( .B1(n174), .B2(n178), .A(n33), .ZN(n958) );
  NAND3_X1 U164 ( .A1(n175), .A2(n179), .A3(warp_id_in[3]), .ZN(n178) );
  OAI21_X1 U165 ( .B1(n167), .B2(n180), .A(n34), .ZN(n957) );
  OAI21_X1 U166 ( .B1(n168), .B2(n180), .A(n35), .ZN(n956) );
  OAI21_X1 U167 ( .B1(n169), .B2(n180), .A(n36), .ZN(n955) );
  OAI21_X1 U168 ( .B1(n170), .B2(n180), .A(n37), .ZN(n954) );
  OAI21_X1 U169 ( .B1(n171), .B2(n180), .A(n38), .ZN(n953) );
  OAI21_X1 U170 ( .B1(n172), .B2(n180), .A(n39), .ZN(n952) );
  OAI21_X1 U171 ( .B1(n173), .B2(n180), .A(n40), .ZN(n951) );
  OAI21_X1 U172 ( .B1(n174), .B2(n180), .A(n41), .ZN(n950) );
  NAND3_X1 U173 ( .A1(n177), .A2(n179), .A3(n175), .ZN(n180) );
  AND4_X1 U174 ( .A1(warp_state_in[0]), .A2(n181), .A3(warp_state_in[1]), .A4(
        n182), .ZN(n175) );
  MUX2_X1 U175 ( .A(warp_checker_state_machine[2]), .B(n183), .S(n145), .Z(
        n1267) );
  OAI221_X1 U176 ( .B1(N567), .B2(n146), .C1(n184), .C2(n185), .A(n186), .ZN(
        n183) );
  OAI221_X1 U177 ( .B1(n7), .B2(n145), .C1(n146), .C2(n147), .A(n187), .ZN(
        n1266) );
  INV_X1 U178 ( .A(N567), .ZN(n147) );
  NAND4_X1 U179 ( .A1(n102), .A2(n187), .A3(n146), .A4(n188), .ZN(n145) );
  AOI21_X1 U180 ( .B1(\warp_cntr[5] ), .B2(n189), .A(n190), .ZN(n188) );
  NAND3_X1 U181 ( .A1(n3), .A2(n8), .A3(warp_checker_state_machine[1]), .ZN(
        n146) );
  OAI21_X1 U182 ( .B1(n988), .B2(n96), .A(n191), .ZN(n1265) );
  NAND2_X1 U183 ( .A1(N703), .A2(n165), .ZN(n191) );
  OAI21_X1 U184 ( .B1(n989), .B2(n96), .A(n192), .ZN(n1264) );
  NAND2_X1 U185 ( .A1(n989), .A2(n165), .ZN(n192) );
  OAI21_X1 U186 ( .B1(n987), .B2(n96), .A(n193), .ZN(n1263) );
  NAND2_X1 U187 ( .A1(N704), .A2(n165), .ZN(n193) );
  OAI21_X1 U188 ( .B1(n986), .B2(n96), .A(n194), .ZN(n1262) );
  NAND2_X1 U189 ( .A1(N705), .A2(n165), .ZN(n194) );
  OAI21_X1 U190 ( .B1(n985), .B2(n96), .A(n195), .ZN(n1261) );
  NAND2_X1 U191 ( .A1(N706), .A2(n165), .ZN(n195) );
  MUX2_X1 U192 ( .A(warp_id_in[0]), .B(warp_id_addr[0]), .S(n101), .Z(n1260)
         );
  MUX2_X1 U193 ( .A(warp_id_in[4]), .B(warp_id_addr[4]), .S(n101), .Z(n1259)
         );
  MUX2_X1 U194 ( .A(warp_id_in[3]), .B(warp_id_addr[3]), .S(n101), .Z(n1258)
         );
  MUX2_X1 U195 ( .A(warp_id_in[2]), .B(warp_id_addr[2]), .S(n101), .Z(n1257)
         );
  MUX2_X1 U196 ( .A(warp_id_in[1]), .B(warp_id_addr[1]), .S(n101), .Z(n1256)
         );
  NAND2_X1 U197 ( .A1(n185), .A2(n196), .ZN(n1255) );
  NAND3_X1 U198 ( .A1(n197), .A2(n102), .A3(pipeline_stall_out), .ZN(n196) );
  INV_X1 U199 ( .A(n181), .ZN(n185) );
  MUX2_X1 U200 ( .A(n96), .B(fence_regs_fence_en_ld[0]), .S(n198), .Z(n1254)
         );
  AOI21_X1 U201 ( .B1(n199), .B2(n200), .A(n201), .ZN(n198) );
  MUX2_X1 U202 ( .A(n96), .B(fence_regs_fence_en_ld[1]), .S(n202), .Z(n1253)
         );
  AOI21_X1 U203 ( .B1(n203), .B2(n200), .A(n204), .ZN(n202) );
  MUX2_X1 U204 ( .A(n96), .B(fence_regs_fence_en_ld[2]), .S(n205), .Z(n1252)
         );
  AOI21_X1 U205 ( .B1(n206), .B2(n200), .A(n207), .ZN(n205) );
  MUX2_X1 U206 ( .A(n96), .B(fence_regs_fence_en_ld[3]), .S(n208), .Z(n1251)
         );
  AOI21_X1 U207 ( .B1(n209), .B2(n200), .A(n210), .ZN(n208) );
  MUX2_X1 U208 ( .A(n96), .B(fence_regs_fence_en_ld[4]), .S(n211), .Z(n1250)
         );
  AOI21_X1 U209 ( .B1(n212), .B2(n200), .A(n213), .ZN(n211) );
  MUX2_X1 U210 ( .A(n96), .B(fence_regs_fence_en_ld[5]), .S(n214), .Z(n1249)
         );
  AOI21_X1 U211 ( .B1(n215), .B2(n200), .A(n216), .ZN(n214) );
  MUX2_X1 U212 ( .A(n96), .B(fence_regs_fence_en_ld[6]), .S(n217), .Z(n1248)
         );
  AOI21_X1 U213 ( .B1(n218), .B2(n200), .A(n219), .ZN(n217) );
  MUX2_X1 U214 ( .A(n96), .B(fence_regs_fence_en_ld[7]), .S(n220), .Z(n1247)
         );
  AOI21_X1 U215 ( .B1(n221), .B2(n200), .A(n222), .ZN(n220) );
  MUX2_X1 U216 ( .A(n97), .B(fence_regs_fence_en_ld[8]), .S(n223), .Z(n1246)
         );
  AOI21_X1 U217 ( .B1(n224), .B2(n199), .A(n225), .ZN(n223) );
  MUX2_X1 U218 ( .A(n97), .B(fence_regs_fence_en_ld[9]), .S(n226), .Z(n1245)
         );
  AOI21_X1 U219 ( .B1(n224), .B2(n203), .A(n227), .ZN(n226) );
  MUX2_X1 U220 ( .A(n97), .B(fence_regs_fence_en_ld[10]), .S(n228), .Z(n1244)
         );
  AOI21_X1 U221 ( .B1(n224), .B2(n206), .A(n229), .ZN(n228) );
  MUX2_X1 U222 ( .A(n97), .B(fence_regs_fence_en_ld[11]), .S(n230), .Z(n1243)
         );
  AOI21_X1 U223 ( .B1(n224), .B2(n209), .A(n231), .ZN(n230) );
  MUX2_X1 U224 ( .A(n97), .B(fence_regs_fence_en_ld[12]), .S(n232), .Z(n1242)
         );
  AOI21_X1 U225 ( .B1(n224), .B2(n212), .A(n233), .ZN(n232) );
  MUX2_X1 U226 ( .A(n97), .B(fence_regs_fence_en_ld[13]), .S(n234), .Z(n1241)
         );
  AOI21_X1 U227 ( .B1(n224), .B2(n215), .A(n235), .ZN(n234) );
  MUX2_X1 U228 ( .A(n97), .B(fence_regs_fence_en_ld[14]), .S(n236), .Z(n1240)
         );
  AOI21_X1 U229 ( .B1(n224), .B2(n218), .A(n237), .ZN(n236) );
  MUX2_X1 U230 ( .A(n97), .B(fence_regs_fence_en_ld[15]), .S(n238), .Z(n1239)
         );
  AOI21_X1 U231 ( .B1(n224), .B2(n221), .A(n239), .ZN(n238) );
  MUX2_X1 U232 ( .A(n97), .B(fence_regs_fence_en_ld[16]), .S(n240), .Z(n1238)
         );
  AOI21_X1 U233 ( .B1(n241), .B2(n199), .A(n242), .ZN(n240) );
  MUX2_X1 U234 ( .A(n97), .B(fence_regs_fence_en_ld[17]), .S(n243), .Z(n1237)
         );
  AOI21_X1 U235 ( .B1(n241), .B2(n203), .A(n244), .ZN(n243) );
  MUX2_X1 U236 ( .A(n97), .B(fence_regs_fence_en_ld[18]), .S(n245), .Z(n1236)
         );
  AOI21_X1 U237 ( .B1(n241), .B2(n206), .A(n246), .ZN(n245) );
  MUX2_X1 U238 ( .A(n97), .B(fence_regs_fence_en_ld[19]), .S(n247), .Z(n1235)
         );
  AOI21_X1 U239 ( .B1(n241), .B2(n209), .A(n248), .ZN(n247) );
  MUX2_X1 U240 ( .A(n97), .B(fence_regs_fence_en_ld[20]), .S(n249), .Z(n1234)
         );
  AOI21_X1 U241 ( .B1(n241), .B2(n212), .A(n250), .ZN(n249) );
  MUX2_X1 U242 ( .A(n97), .B(fence_regs_fence_en_ld[21]), .S(n251), .Z(n1233)
         );
  AOI21_X1 U243 ( .B1(n241), .B2(n215), .A(n252), .ZN(n251) );
  MUX2_X1 U244 ( .A(n97), .B(fence_regs_fence_en_ld[22]), .S(n253), .Z(n1232)
         );
  AOI21_X1 U245 ( .B1(n241), .B2(n218), .A(n254), .ZN(n253) );
  MUX2_X1 U246 ( .A(n97), .B(fence_regs_fence_en_ld[23]), .S(n255), .Z(n1231)
         );
  AOI21_X1 U247 ( .B1(n241), .B2(n221), .A(n256), .ZN(n255) );
  AND3_X1 U248 ( .A1(warp_id_addr[4]), .A2(n6), .A3(n257), .ZN(n241) );
  MUX2_X1 U249 ( .A(n98), .B(fence_regs_fence_en_ld[24]), .S(n258), .Z(n1230)
         );
  AOI21_X1 U250 ( .B1(n259), .B2(n199), .A(n260), .ZN(n258) );
  NOR3_X1 U251 ( .A1(warp_id_addr[1]), .A2(warp_id_addr[2]), .A3(
        warp_id_addr[0]), .ZN(n199) );
  MUX2_X1 U252 ( .A(n98), .B(fence_regs_fence_en_ld[25]), .S(n261), .Z(n1229)
         );
  AOI21_X1 U253 ( .B1(n259), .B2(n203), .A(n262), .ZN(n261) );
  NOR3_X1 U254 ( .A1(warp_id_addr[1]), .A2(warp_id_addr[2]), .A3(n4), .ZN(n203) );
  MUX2_X1 U255 ( .A(n98), .B(fence_regs_fence_en_ld[26]), .S(n263), .Z(n1228)
         );
  AOI21_X1 U256 ( .B1(n259), .B2(n206), .A(n264), .ZN(n263) );
  NOR3_X1 U257 ( .A1(warp_id_addr[0]), .A2(warp_id_addr[2]), .A3(n5), .ZN(n206) );
  MUX2_X1 U258 ( .A(n98), .B(fence_regs_fence_en_ld[27]), .S(n265), .Z(n1227)
         );
  AOI21_X1 U259 ( .B1(n259), .B2(n209), .A(n266), .ZN(n265) );
  NOR3_X1 U260 ( .A1(n4), .A2(warp_id_addr[2]), .A3(n5), .ZN(n209) );
  MUX2_X1 U261 ( .A(n98), .B(fence_regs_fence_en_ld[28]), .S(n267), .Z(n1226)
         );
  AOI21_X1 U262 ( .B1(n259), .B2(n212), .A(n268), .ZN(n267) );
  AND3_X1 U263 ( .A1(n4), .A2(n5), .A3(warp_id_addr[2]), .ZN(n212) );
  MUX2_X1 U264 ( .A(n98), .B(fence_regs_fence_en_ld[29]), .S(n269), .Z(n1225)
         );
  AOI21_X1 U265 ( .B1(n259), .B2(n215), .A(n270), .ZN(n269) );
  AND3_X1 U266 ( .A1(warp_id_addr[0]), .A2(n5), .A3(warp_id_addr[2]), .ZN(n215) );
  MUX2_X1 U267 ( .A(n98), .B(fence_regs_fence_en_ld[30]), .S(n271), .Z(n1224)
         );
  AOI21_X1 U268 ( .B1(n259), .B2(n218), .A(n272), .ZN(n271) );
  AND3_X1 U269 ( .A1(warp_id_addr[2]), .A2(n4), .A3(warp_id_addr[1]), .ZN(n218) );
  MUX2_X1 U270 ( .A(n98), .B(fence_regs_fence_en_ld[31]), .S(n273), .Z(n1223)
         );
  AOI21_X1 U271 ( .B1(n259), .B2(n221), .A(n274), .ZN(n273) );
  AND3_X1 U272 ( .A1(warp_id_addr[2]), .A2(warp_id_addr[0]), .A3(
        warp_id_addr[1]), .ZN(n221) );
  AND3_X1 U273 ( .A1(warp_id_addr[3]), .A2(warp_id_addr[4]), .A3(n257), .ZN(
        n259) );
  NAND2_X1 U274 ( .A1(n186), .A2(n102), .ZN(n163) );
  INV_X1 U275 ( .A(n189), .ZN(n186) );
  OAI22_X1 U276 ( .A1(n78), .A2(n781), .B1(n84), .B2(n275), .ZN(n1222) );
  OAI22_X1 U277 ( .A1(n77), .A2(n782), .B1(n83), .B2(n144), .ZN(n1221) );
  OAI22_X1 U278 ( .A1(n77), .A2(n783), .B1(n84), .B2(n142), .ZN(n1220) );
  OAI22_X1 U279 ( .A1(n77), .A2(n784), .B1(n84), .B2(n140), .ZN(n1219) );
  OAI22_X1 U280 ( .A1(n77), .A2(n785), .B1(n84), .B2(n138), .ZN(n1218) );
  OAI22_X1 U281 ( .A1(n77), .A2(n786), .B1(n84), .B2(n276), .ZN(n1217) );
  OAI21_X1 U282 ( .B1(n82), .B2(n787), .A(n83), .ZN(n1216) );
  OAI22_X1 U283 ( .A1(n77), .A2(n788), .B1(n84), .B2(n179), .ZN(n1215) );
  OAI22_X1 U284 ( .A1(n77), .A2(n789), .B1(n84), .B2(n177), .ZN(n1214) );
  OAI22_X1 U285 ( .A1(n77), .A2(n790), .B1(n84), .B2(n277), .ZN(n1213) );
  OAI222_X1 U286 ( .A1(n989), .A2(n278), .B1(n162), .B2(n275), .C1(n160), .C2(
        n791), .ZN(n1212) );
  OAI21_X1 U287 ( .B1(n160), .B2(n1173), .A(n279), .ZN(n1211) );
  NAND3_X1 U288 ( .A1(n280), .A2(warp_state_in[1]), .A3(warp_state_in[0]), 
        .ZN(n279) );
  INV_X1 U289 ( .A(n162), .ZN(n280) );
  OAI222_X1 U290 ( .A1(n985), .A2(n278), .B1(n162), .B2(n179), .C1(n160), .C2(
        n792), .ZN(n1210) );
  OAI222_X1 U291 ( .A1(n986), .A2(n278), .B1(n162), .B2(n177), .C1(n160), .C2(
        n793), .ZN(n1209) );
  OAI222_X1 U292 ( .A1(n987), .A2(n278), .B1(n162), .B2(n277), .C1(n160), .C2(
        n794), .ZN(n1208) );
  OAI222_X1 U293 ( .A1(n988), .A2(n278), .B1(n162), .B2(n276), .C1(n160), .C2(
        n795), .ZN(n1207) );
  NAND2_X1 U294 ( .A1(n181), .A2(n160), .ZN(n162) );
  NAND2_X1 U295 ( .A1(n189), .A2(n160), .ZN(n278) );
  OAI211_X1 U296 ( .C1(n796), .C2(n282), .A(n281), .B(n83), .ZN(n1206) );
  NAND2_X1 U297 ( .A1(n1), .A2(n283), .ZN(n282) );
  MUX2_X1 U298 ( .A(fence_regs_fence_en_out[0]), .B(n100), .S(n201), .Z(n1205)
         );
  OAI22_X1 U299 ( .A1(n174), .A2(n284), .B1(n285), .B2(n286), .ZN(n201) );
  MUX2_X1 U300 ( .A(fence_regs_fence_en_out[31]), .B(n100), .S(n274), .Z(n1204) );
  OAI22_X1 U301 ( .A1(n167), .A2(n287), .B1(n288), .B2(n289), .ZN(n274) );
  MUX2_X1 U302 ( .A(fence_regs_fence_en_out[30]), .B(n100), .S(n272), .Z(n1203) );
  OAI22_X1 U303 ( .A1(n168), .A2(n287), .B1(n290), .B2(n289), .ZN(n272) );
  MUX2_X1 U304 ( .A(fence_regs_fence_en_out[29]), .B(n100), .S(n270), .Z(n1202) );
  OAI22_X1 U305 ( .A1(n169), .A2(n287), .B1(n291), .B2(n289), .ZN(n270) );
  MUX2_X1 U306 ( .A(fence_regs_fence_en_out[28]), .B(n100), .S(n268), .Z(n1201) );
  OAI22_X1 U307 ( .A1(n170), .A2(n287), .B1(n292), .B2(n289), .ZN(n268) );
  MUX2_X1 U308 ( .A(fence_regs_fence_en_out[27]), .B(n100), .S(n266), .Z(n1200) );
  OAI22_X1 U309 ( .A1(n171), .A2(n287), .B1(n293), .B2(n289), .ZN(n266) );
  MUX2_X1 U310 ( .A(fence_regs_fence_en_out[26]), .B(n100), .S(n264), .Z(n1199) );
  OAI22_X1 U311 ( .A1(n172), .A2(n287), .B1(n294), .B2(n289), .ZN(n264) );
  MUX2_X1 U312 ( .A(fence_regs_fence_en_out[25]), .B(n100), .S(n262), .Z(n1198) );
  OAI22_X1 U313 ( .A1(n173), .A2(n287), .B1(n295), .B2(n289), .ZN(n262) );
  MUX2_X1 U314 ( .A(fence_regs_fence_en_out[24]), .B(n100), .S(n260), .Z(n1197) );
  OAI22_X1 U315 ( .A1(n174), .A2(n287), .B1(n285), .B2(n289), .ZN(n260) );
  NAND3_X1 U316 ( .A1(N116), .A2(N115), .A3(n296), .ZN(n289) );
  NAND3_X1 U317 ( .A1(warp_id_in[4]), .A2(warp_id_in[3]), .A3(n297), .ZN(n287)
         );
  MUX2_X1 U318 ( .A(fence_regs_fence_en_out[23]), .B(n100), .S(n256), .Z(n1196) );
  OAI22_X1 U319 ( .A1(n167), .A2(n298), .B1(n288), .B2(n299), .ZN(n256) );
  MUX2_X1 U320 ( .A(fence_regs_fence_en_out[22]), .B(n100), .S(n254), .Z(n1195) );
  OAI22_X1 U321 ( .A1(n168), .A2(n298), .B1(n290), .B2(n299), .ZN(n254) );
  MUX2_X1 U322 ( .A(fence_regs_fence_en_out[21]), .B(n100), .S(n252), .Z(n1194) );
  OAI22_X1 U323 ( .A1(n169), .A2(n298), .B1(n291), .B2(n299), .ZN(n252) );
  MUX2_X1 U324 ( .A(fence_regs_fence_en_out[20]), .B(n100), .S(n250), .Z(n1193) );
  OAI22_X1 U325 ( .A1(n170), .A2(n298), .B1(n292), .B2(n299), .ZN(n250) );
  MUX2_X1 U326 ( .A(fence_regs_fence_en_out[19]), .B(n100), .S(n248), .Z(n1192) );
  OAI22_X1 U327 ( .A1(n171), .A2(n298), .B1(n293), .B2(n299), .ZN(n248) );
  MUX2_X1 U328 ( .A(fence_regs_fence_en_out[18]), .B(n100), .S(n246), .Z(n1191) );
  OAI22_X1 U329 ( .A1(n172), .A2(n298), .B1(n294), .B2(n299), .ZN(n246) );
  MUX2_X1 U330 ( .A(fence_regs_fence_en_out[17]), .B(n100), .S(n244), .Z(n1190) );
  OAI22_X1 U331 ( .A1(n173), .A2(n298), .B1(n295), .B2(n299), .ZN(n244) );
  MUX2_X1 U332 ( .A(fence_regs_fence_en_out[16]), .B(n100), .S(n242), .Z(n1189) );
  OAI22_X1 U333 ( .A1(n174), .A2(n298), .B1(n285), .B2(n299), .ZN(n242) );
  NAND3_X1 U334 ( .A1(n296), .A2(N116), .A3(n986), .ZN(n299) );
  NAND3_X1 U335 ( .A1(warp_id_in[4]), .A2(n177), .A3(n297), .ZN(n298) );
  MUX2_X1 U336 ( .A(fence_regs_fence_en_out[15]), .B(n100), .S(n239), .Z(n1188) );
  OAI22_X1 U337 ( .A1(n167), .A2(n300), .B1(n288), .B2(n301), .ZN(n239) );
  MUX2_X1 U338 ( .A(fence_regs_fence_en_out[14]), .B(n99), .S(n237), .Z(n1187)
         );
  OAI22_X1 U339 ( .A1(n168), .A2(n300), .B1(n290), .B2(n301), .ZN(n237) );
  MUX2_X1 U340 ( .A(fence_regs_fence_en_out[13]), .B(n99), .S(n235), .Z(n1186)
         );
  OAI22_X1 U341 ( .A1(n169), .A2(n300), .B1(n291), .B2(n301), .ZN(n235) );
  MUX2_X1 U342 ( .A(fence_regs_fence_en_out[12]), .B(n99), .S(n233), .Z(n1185)
         );
  OAI22_X1 U343 ( .A1(n170), .A2(n300), .B1(n292), .B2(n301), .ZN(n233) );
  MUX2_X1 U344 ( .A(fence_regs_fence_en_out[11]), .B(n99), .S(n231), .Z(n1184)
         );
  OAI22_X1 U345 ( .A1(n171), .A2(n300), .B1(n293), .B2(n301), .ZN(n231) );
  MUX2_X1 U346 ( .A(fence_regs_fence_en_out[10]), .B(n99), .S(n229), .Z(n1183)
         );
  OAI22_X1 U347 ( .A1(n172), .A2(n300), .B1(n294), .B2(n301), .ZN(n229) );
  MUX2_X1 U348 ( .A(fence_regs_fence_en_out[9]), .B(n99), .S(n227), .Z(n1182)
         );
  OAI22_X1 U349 ( .A1(n173), .A2(n300), .B1(n295), .B2(n301), .ZN(n227) );
  MUX2_X1 U350 ( .A(fence_regs_fence_en_out[8]), .B(n99), .S(n225), .Z(n1181)
         );
  OAI22_X1 U351 ( .A1(n174), .A2(n300), .B1(n285), .B2(n301), .ZN(n225) );
  NAND3_X1 U352 ( .A1(n296), .A2(N115), .A3(n985), .ZN(n301) );
  NAND3_X1 U353 ( .A1(n988), .A2(n987), .A3(n989), .ZN(n285) );
  NAND3_X1 U354 ( .A1(warp_id_in[3]), .A2(n179), .A3(n297), .ZN(n300) );
  NAND3_X1 U355 ( .A1(n276), .A2(n277), .A3(n275), .ZN(n174) );
  MUX2_X1 U356 ( .A(fence_regs_fence_en_out[7]), .B(n99), .S(n222), .Z(n1180)
         );
  OAI22_X1 U357 ( .A1(n167), .A2(n284), .B1(n286), .B2(n288), .ZN(n222) );
  NAND3_X1 U358 ( .A1(N113), .A2(N112), .A3(N114), .ZN(n288) );
  NAND3_X1 U359 ( .A1(warp_id_in[1]), .A2(warp_id_in[0]), .A3(warp_id_in[2]), 
        .ZN(n167) );
  MUX2_X1 U360 ( .A(fence_regs_fence_en_out[6]), .B(n99), .S(n219), .Z(n1179)
         );
  OAI22_X1 U361 ( .A1(n168), .A2(n284), .B1(n286), .B2(n290), .ZN(n219) );
  NAND3_X1 U362 ( .A1(N114), .A2(N113), .A3(n989), .ZN(n290) );
  NAND3_X1 U363 ( .A1(warp_id_in[1]), .A2(n275), .A3(warp_id_in[2]), .ZN(n168)
         );
  MUX2_X1 U364 ( .A(fence_regs_fence_en_out[5]), .B(n99), .S(n216), .Z(n1178)
         );
  OAI22_X1 U365 ( .A1(n169), .A2(n284), .B1(n286), .B2(n291), .ZN(n216) );
  NAND3_X1 U366 ( .A1(N114), .A2(N112), .A3(n988), .ZN(n291) );
  NAND3_X1 U367 ( .A1(warp_id_in[0]), .A2(n276), .A3(warp_id_in[2]), .ZN(n169)
         );
  MUX2_X1 U368 ( .A(fence_regs_fence_en_out[4]), .B(n99), .S(n213), .Z(n1177)
         );
  OAI22_X1 U369 ( .A1(n170), .A2(n284), .B1(n286), .B2(n292), .ZN(n213) );
  NAND3_X1 U370 ( .A1(n988), .A2(N114), .A3(n989), .ZN(n292) );
  NAND3_X1 U371 ( .A1(n275), .A2(n276), .A3(warp_id_in[2]), .ZN(n170) );
  MUX2_X1 U372 ( .A(fence_regs_fence_en_out[3]), .B(n99), .S(n210), .Z(n1176)
         );
  OAI22_X1 U373 ( .A1(n171), .A2(n284), .B1(n286), .B2(n293), .ZN(n210) );
  NAND3_X1 U374 ( .A1(N113), .A2(N112), .A3(n987), .ZN(n293) );
  NAND3_X1 U375 ( .A1(warp_id_in[0]), .A2(n277), .A3(warp_id_in[1]), .ZN(n171)
         );
  MUX2_X1 U376 ( .A(fence_regs_fence_en_out[2]), .B(n99), .S(n207), .Z(n1175)
         );
  OAI22_X1 U377 ( .A1(n172), .A2(n284), .B1(n286), .B2(n294), .ZN(n207) );
  NAND3_X1 U378 ( .A1(n987), .A2(N113), .A3(n989), .ZN(n294) );
  NAND3_X1 U379 ( .A1(n275), .A2(n277), .A3(warp_id_in[1]), .ZN(n172) );
  INV_X1 U380 ( .A(warp_id_in[0]), .ZN(n275) );
  MUX2_X1 U381 ( .A(fence_regs_fence_en_out[1]), .B(n99), .S(n204), .Z(n1174)
         );
  OAI22_X1 U382 ( .A1(n173), .A2(n284), .B1(n286), .B2(n295), .ZN(n204) );
  NAND3_X1 U383 ( .A1(n987), .A2(N112), .A3(n988), .ZN(n295) );
  NAND3_X1 U384 ( .A1(n985), .A2(n296), .A3(n986), .ZN(n286) );
  INV_X1 U385 ( .A(n281), .ZN(n296) );
  NAND2_X1 U386 ( .A1(N572), .A2(n165), .ZN(n281) );
  INV_X1 U387 ( .A(n283), .ZN(n165) );
  NAND2_X1 U388 ( .A1(n9), .A2(n189), .ZN(n283) );
  NOR3_X1 U389 ( .A1(n3), .A2(warp_checker_state_machine[2]), .A3(n7), .ZN(
        n189) );
  NAND3_X1 U390 ( .A1(n177), .A2(n179), .A3(n297), .ZN(n284) );
  INV_X1 U391 ( .A(n148), .ZN(n297) );
  NAND2_X1 U392 ( .A1(n181), .A2(n184), .ZN(n148) );
  NOR3_X1 U393 ( .A1(n302), .A2(warp_state_in[0]), .A3(n161), .ZN(n184) );
  INV_X1 U394 ( .A(warp_state_in[1]), .ZN(n161) );
  INV_X1 U395 ( .A(warp_id_in[4]), .ZN(n179) );
  INV_X1 U396 ( .A(warp_id_in[3]), .ZN(n177) );
  NAND3_X1 U397 ( .A1(n276), .A2(n277), .A3(warp_id_in[0]), .ZN(n173) );
  INV_X1 U398 ( .A(warp_id_in[2]), .ZN(n277) );
  INV_X1 U399 ( .A(warp_id_in[1]), .ZN(n276) );
  MUX2_X1 U400 ( .A(warps_done_mask[0]), .B(warps_done_mask_out[0]), .S(n106), 
        .Z(n1140) );
  MUX2_X1 U401 ( .A(warps_done_mask[1]), .B(warps_done_mask_out[1]), .S(n106), 
        .Z(n1139) );
  MUX2_X1 U402 ( .A(warps_done_mask[2]), .B(warps_done_mask_out[2]), .S(n106), 
        .Z(n1138) );
  MUX2_X1 U403 ( .A(warps_done_mask[3]), .B(warps_done_mask_out[3]), .S(n106), 
        .Z(n1137) );
  MUX2_X1 U404 ( .A(warps_done_mask[4]), .B(warps_done_mask_out[4]), .S(n106), 
        .Z(n1136) );
  MUX2_X1 U405 ( .A(warps_done_mask[5]), .B(warps_done_mask_out[5]), .S(n106), 
        .Z(n1135) );
  MUX2_X1 U406 ( .A(warps_done_mask[6]), .B(warps_done_mask_out[6]), .S(n106), 
        .Z(n1134) );
  MUX2_X1 U407 ( .A(warps_done_mask[7]), .B(warps_done_mask_out[7]), .S(n106), 
        .Z(n1133) );
  MUX2_X1 U408 ( .A(warps_done_mask[8]), .B(warps_done_mask_out[8]), .S(n105), 
        .Z(n1132) );
  MUX2_X1 U409 ( .A(warps_done_mask[9]), .B(warps_done_mask_out[9]), .S(n105), 
        .Z(n1131) );
  MUX2_X1 U410 ( .A(warps_done_mask[10]), .B(warps_done_mask_out[10]), .S(n105), .Z(n1130) );
  MUX2_X1 U411 ( .A(warps_done_mask[11]), .B(warps_done_mask_out[11]), .S(n105), .Z(n1129) );
  MUX2_X1 U412 ( .A(warps_done_mask[12]), .B(warps_done_mask_out[12]), .S(n105), .Z(n1128) );
  MUX2_X1 U413 ( .A(warps_done_mask[13]), .B(warps_done_mask_out[13]), .S(n105), .Z(n1127) );
  MUX2_X1 U414 ( .A(warps_done_mask[14]), .B(warps_done_mask_out[14]), .S(n105), .Z(n1126) );
  MUX2_X1 U415 ( .A(warps_done_mask[15]), .B(warps_done_mask_out[15]), .S(n105), .Z(n1125) );
  MUX2_X1 U416 ( .A(warps_done_mask[16]), .B(warps_done_mask_out[16]), .S(n105), .Z(n1124) );
  MUX2_X1 U417 ( .A(warps_done_mask[17]), .B(warps_done_mask_out[17]), .S(n105), .Z(n1123) );
  MUX2_X1 U418 ( .A(warps_done_mask[18]), .B(warps_done_mask_out[18]), .S(n105), .Z(n1122) );
  MUX2_X1 U419 ( .A(warps_done_mask[19]), .B(warps_done_mask_out[19]), .S(n105), .Z(n1121) );
  MUX2_X1 U420 ( .A(warps_done_mask[20]), .B(warps_done_mask_out[20]), .S(n104), .Z(n1120) );
  MUX2_X1 U421 ( .A(warps_done_mask[21]), .B(warps_done_mask_out[21]), .S(n104), .Z(n1119) );
  MUX2_X1 U422 ( .A(warps_done_mask[22]), .B(warps_done_mask_out[22]), .S(n104), .Z(n1118) );
  MUX2_X1 U423 ( .A(warps_done_mask[23]), .B(warps_done_mask_out[23]), .S(n104), .Z(n1117) );
  MUX2_X1 U424 ( .A(warps_done_mask[24]), .B(warps_done_mask_out[24]), .S(n104), .Z(n1116) );
  MUX2_X1 U425 ( .A(warps_done_mask[25]), .B(warps_done_mask_out[25]), .S(n104), .Z(n1115) );
  MUX2_X1 U426 ( .A(warps_done_mask[26]), .B(warps_done_mask_out[26]), .S(n104), .Z(n1114) );
  MUX2_X1 U427 ( .A(warps_done_mask[27]), .B(warps_done_mask_out[27]), .S(n104), .Z(n1113) );
  MUX2_X1 U428 ( .A(warps_done_mask[28]), .B(warps_done_mask_out[28]), .S(n104), .Z(n1112) );
  MUX2_X1 U429 ( .A(warps_done_mask[29]), .B(warps_done_mask_out[29]), .S(n104), .Z(n1111) );
  MUX2_X1 U430 ( .A(warps_done_mask[30]), .B(warps_done_mask_out[30]), .S(n104), .Z(n1110) );
  MUX2_X1 U431 ( .A(warps_done_mask[31]), .B(warps_done_mask_out[31]), .S(n104), .Z(n1109) );
  AOI21_X1 U432 ( .B1(n304), .B2(n99), .A(n190), .ZN(n303) );
  OAI22_X1 U433 ( .A1(n77), .A2(n916), .B1(n84), .B2(n305), .ZN(n1108) );
  INV_X1 U434 ( .A(current_mask_in[0]), .ZN(n305) );
  OAI22_X1 U435 ( .A1(n77), .A2(n915), .B1(n84), .B2(n306), .ZN(n1107) );
  INV_X1 U436 ( .A(current_mask_in[1]), .ZN(n306) );
  OAI22_X1 U437 ( .A1(n77), .A2(n914), .B1(n84), .B2(n307), .ZN(n1106) );
  INV_X1 U438 ( .A(current_mask_in[2]), .ZN(n307) );
  OAI22_X1 U439 ( .A1(n77), .A2(n913), .B1(n85), .B2(n308), .ZN(n1105) );
  INV_X1 U440 ( .A(current_mask_in[3]), .ZN(n308) );
  OAI22_X1 U441 ( .A1(n78), .A2(n912), .B1(n85), .B2(n309), .ZN(n1104) );
  INV_X1 U442 ( .A(current_mask_in[4]), .ZN(n309) );
  OAI22_X1 U443 ( .A1(n78), .A2(n911), .B1(n85), .B2(n310), .ZN(n1103) );
  INV_X1 U444 ( .A(current_mask_in[5]), .ZN(n310) );
  OAI22_X1 U445 ( .A1(n78), .A2(n910), .B1(n85), .B2(n311), .ZN(n1102) );
  INV_X1 U446 ( .A(current_mask_in[6]), .ZN(n311) );
  OAI22_X1 U447 ( .A1(n78), .A2(n909), .B1(n85), .B2(n312), .ZN(n1101) );
  INV_X1 U448 ( .A(current_mask_in[7]), .ZN(n312) );
  OAI22_X1 U449 ( .A1(n78), .A2(n908), .B1(n85), .B2(n313), .ZN(n1100) );
  INV_X1 U450 ( .A(current_mask_in[8]), .ZN(n313) );
  OAI22_X1 U451 ( .A1(n78), .A2(n907), .B1(n85), .B2(n314), .ZN(n1099) );
  INV_X1 U452 ( .A(current_mask_in[9]), .ZN(n314) );
  OAI22_X1 U453 ( .A1(n78), .A2(n906), .B1(n85), .B2(n315), .ZN(n1098) );
  INV_X1 U454 ( .A(current_mask_in[10]), .ZN(n315) );
  OAI22_X1 U455 ( .A1(n78), .A2(n905), .B1(n85), .B2(n316), .ZN(n1097) );
  INV_X1 U456 ( .A(current_mask_in[11]), .ZN(n316) );
  OAI22_X1 U457 ( .A1(n78), .A2(n904), .B1(n85), .B2(n317), .ZN(n1096) );
  INV_X1 U458 ( .A(current_mask_in[12]), .ZN(n317) );
  OAI22_X1 U459 ( .A1(n78), .A2(n903), .B1(n85), .B2(n318), .ZN(n1095) );
  INV_X1 U460 ( .A(current_mask_in[13]), .ZN(n318) );
  OAI22_X1 U461 ( .A1(n78), .A2(n902), .B1(n85), .B2(n319), .ZN(n1094) );
  INV_X1 U462 ( .A(current_mask_in[14]), .ZN(n319) );
  OAI22_X1 U463 ( .A1(n78), .A2(n901), .B1(n86), .B2(n320), .ZN(n1093) );
  INV_X1 U464 ( .A(current_mask_in[15]), .ZN(n320) );
  OAI22_X1 U465 ( .A1(n79), .A2(n900), .B1(n86), .B2(n321), .ZN(n1092) );
  INV_X1 U466 ( .A(current_mask_in[16]), .ZN(n321) );
  OAI22_X1 U467 ( .A1(n79), .A2(n899), .B1(n86), .B2(n322), .ZN(n1091) );
  INV_X1 U468 ( .A(current_mask_in[17]), .ZN(n322) );
  OAI22_X1 U469 ( .A1(n79), .A2(n898), .B1(n86), .B2(n323), .ZN(n1090) );
  INV_X1 U470 ( .A(current_mask_in[18]), .ZN(n323) );
  OAI22_X1 U471 ( .A1(n79), .A2(n897), .B1(n86), .B2(n324), .ZN(n1089) );
  INV_X1 U472 ( .A(current_mask_in[19]), .ZN(n324) );
  OAI22_X1 U473 ( .A1(n79), .A2(n896), .B1(n86), .B2(n325), .ZN(n1088) );
  INV_X1 U474 ( .A(current_mask_in[20]), .ZN(n325) );
  OAI22_X1 U475 ( .A1(n79), .A2(n895), .B1(n86), .B2(n326), .ZN(n1087) );
  INV_X1 U476 ( .A(current_mask_in[21]), .ZN(n326) );
  OAI22_X1 U477 ( .A1(n79), .A2(n894), .B1(n86), .B2(n327), .ZN(n1086) );
  INV_X1 U478 ( .A(current_mask_in[22]), .ZN(n327) );
  OAI22_X1 U479 ( .A1(n79), .A2(n893), .B1(n86), .B2(n328), .ZN(n1085) );
  INV_X1 U480 ( .A(current_mask_in[23]), .ZN(n328) );
  OAI22_X1 U481 ( .A1(n79), .A2(n892), .B1(n86), .B2(n329), .ZN(n1084) );
  INV_X1 U482 ( .A(current_mask_in[24]), .ZN(n329) );
  OAI22_X1 U483 ( .A1(n79), .A2(n891), .B1(n86), .B2(n330), .ZN(n1083) );
  INV_X1 U484 ( .A(current_mask_in[25]), .ZN(n330) );
  OAI22_X1 U485 ( .A1(n79), .A2(n890), .B1(n86), .B2(n331), .ZN(n1082) );
  INV_X1 U486 ( .A(current_mask_in[26]), .ZN(n331) );
  OAI22_X1 U487 ( .A1(n79), .A2(n889), .B1(n87), .B2(n332), .ZN(n1081) );
  INV_X1 U488 ( .A(current_mask_in[27]), .ZN(n332) );
  OAI22_X1 U489 ( .A1(n79), .A2(n888), .B1(n87), .B2(n333), .ZN(n1080) );
  INV_X1 U490 ( .A(current_mask_in[28]), .ZN(n333) );
  OAI22_X1 U491 ( .A1(n82), .A2(n887), .B1(n87), .B2(n334), .ZN(n1079) );
  INV_X1 U492 ( .A(current_mask_in[29]), .ZN(n334) );
  OAI22_X1 U493 ( .A1(n81), .A2(n886), .B1(n87), .B2(n335), .ZN(n1078) );
  INV_X1 U494 ( .A(current_mask_in[30]), .ZN(n335) );
  OAI22_X1 U495 ( .A1(n80), .A2(n885), .B1(n87), .B2(n336), .ZN(n1077) );
  INV_X1 U496 ( .A(current_mask_in[31]), .ZN(n336) );
  OAI22_X1 U497 ( .A1(n78), .A2(n884), .B1(n87), .B2(n337), .ZN(n1076) );
  INV_X1 U498 ( .A(initial_mask_in[0]), .ZN(n337) );
  OAI22_X1 U499 ( .A1(n77), .A2(n883), .B1(n87), .B2(n338), .ZN(n1075) );
  INV_X1 U500 ( .A(initial_mask_in[1]), .ZN(n338) );
  OAI22_X1 U501 ( .A1(n79), .A2(n882), .B1(n87), .B2(n339), .ZN(n1074) );
  INV_X1 U502 ( .A(initial_mask_in[2]), .ZN(n339) );
  OAI22_X1 U503 ( .A1(n82), .A2(n881), .B1(n87), .B2(n340), .ZN(n1073) );
  INV_X1 U504 ( .A(initial_mask_in[3]), .ZN(n340) );
  OAI22_X1 U505 ( .A1(n81), .A2(n880), .B1(n87), .B2(n341), .ZN(n1072) );
  INV_X1 U506 ( .A(initial_mask_in[4]), .ZN(n341) );
  OAI22_X1 U507 ( .A1(n80), .A2(n879), .B1(n87), .B2(n342), .ZN(n1071) );
  INV_X1 U508 ( .A(initial_mask_in[5]), .ZN(n342) );
  OAI22_X1 U509 ( .A1(n81), .A2(n878), .B1(n87), .B2(n343), .ZN(n1070) );
  INV_X1 U510 ( .A(initial_mask_in[6]), .ZN(n343) );
  OAI22_X1 U511 ( .A1(n80), .A2(n877), .B1(n88), .B2(n344), .ZN(n1069) );
  INV_X1 U512 ( .A(initial_mask_in[7]), .ZN(n344) );
  OAI22_X1 U513 ( .A1(n77), .A2(n876), .B1(n88), .B2(n345), .ZN(n1068) );
  INV_X1 U514 ( .A(initial_mask_in[8]), .ZN(n345) );
  OAI22_X1 U515 ( .A1(n79), .A2(n875), .B1(n88), .B2(n346), .ZN(n1067) );
  INV_X1 U516 ( .A(initial_mask_in[9]), .ZN(n346) );
  OAI22_X1 U517 ( .A1(n81), .A2(n874), .B1(n88), .B2(n347), .ZN(n1066) );
  INV_X1 U518 ( .A(initial_mask_in[10]), .ZN(n347) );
  OAI22_X1 U519 ( .A1(n80), .A2(n873), .B1(n88), .B2(n348), .ZN(n1065) );
  INV_X1 U520 ( .A(initial_mask_in[11]), .ZN(n348) );
  OAI22_X1 U521 ( .A1(n77), .A2(n872), .B1(n88), .B2(n349), .ZN(n1064) );
  INV_X1 U522 ( .A(initial_mask_in[12]), .ZN(n349) );
  OAI22_X1 U523 ( .A1(n78), .A2(n871), .B1(n88), .B2(n350), .ZN(n1063) );
  INV_X1 U524 ( .A(initial_mask_in[13]), .ZN(n350) );
  OAI22_X1 U525 ( .A1(n77), .A2(n870), .B1(n88), .B2(n351), .ZN(n1062) );
  INV_X1 U526 ( .A(initial_mask_in[14]), .ZN(n351) );
  OAI22_X1 U527 ( .A1(n79), .A2(n869), .B1(n88), .B2(n352), .ZN(n1061) );
  INV_X1 U528 ( .A(initial_mask_in[15]), .ZN(n352) );
  OAI22_X1 U529 ( .A1(n81), .A2(n868), .B1(n88), .B2(n353), .ZN(n1060) );
  INV_X1 U530 ( .A(initial_mask_in[16]), .ZN(n353) );
  OAI22_X1 U531 ( .A1(n80), .A2(n867), .B1(n88), .B2(n354), .ZN(n1059) );
  INV_X1 U532 ( .A(initial_mask_in[17]), .ZN(n354) );
  OAI22_X1 U533 ( .A1(n79), .A2(n866), .B1(n89), .B2(n355), .ZN(n1058) );
  INV_X1 U534 ( .A(initial_mask_in[18]), .ZN(n355) );
  OAI22_X1 U535 ( .A1(n80), .A2(n865), .B1(n89), .B2(n356), .ZN(n1057) );
  INV_X1 U536 ( .A(initial_mask_in[19]), .ZN(n356) );
  OAI22_X1 U537 ( .A1(n80), .A2(n864), .B1(n89), .B2(n357), .ZN(n1056) );
  INV_X1 U538 ( .A(initial_mask_in[20]), .ZN(n357) );
  OAI22_X1 U539 ( .A1(n80), .A2(n863), .B1(n89), .B2(n358), .ZN(n1055) );
  INV_X1 U540 ( .A(initial_mask_in[21]), .ZN(n358) );
  OAI22_X1 U541 ( .A1(n80), .A2(n862), .B1(n89), .B2(n359), .ZN(n1054) );
  INV_X1 U542 ( .A(initial_mask_in[22]), .ZN(n359) );
  OAI22_X1 U543 ( .A1(n80), .A2(n861), .B1(n89), .B2(n360), .ZN(n1053) );
  INV_X1 U544 ( .A(initial_mask_in[23]), .ZN(n360) );
  OAI22_X1 U545 ( .A1(n80), .A2(n860), .B1(n89), .B2(n361), .ZN(n1052) );
  INV_X1 U546 ( .A(initial_mask_in[24]), .ZN(n361) );
  OAI22_X1 U547 ( .A1(n80), .A2(n859), .B1(n89), .B2(n362), .ZN(n1051) );
  INV_X1 U548 ( .A(initial_mask_in[25]), .ZN(n362) );
  OAI22_X1 U549 ( .A1(n80), .A2(n858), .B1(n89), .B2(n363), .ZN(n1050) );
  INV_X1 U550 ( .A(initial_mask_in[26]), .ZN(n363) );
  OAI22_X1 U551 ( .A1(n80), .A2(n857), .B1(n89), .B2(n364), .ZN(n1049) );
  INV_X1 U552 ( .A(initial_mask_in[27]), .ZN(n364) );
  OAI22_X1 U553 ( .A1(n80), .A2(n856), .B1(n89), .B2(n365), .ZN(n1048) );
  INV_X1 U554 ( .A(initial_mask_in[28]), .ZN(n365) );
  OAI22_X1 U555 ( .A1(n80), .A2(n855), .B1(n89), .B2(n366), .ZN(n1047) );
  INV_X1 U556 ( .A(initial_mask_in[29]), .ZN(n366) );
  OAI22_X1 U557 ( .A1(n80), .A2(n854), .B1(n90), .B2(n367), .ZN(n1046) );
  INV_X1 U558 ( .A(initial_mask_in[30]), .ZN(n367) );
  OAI22_X1 U559 ( .A1(n81), .A2(n853), .B1(n90), .B2(n368), .ZN(n1045) );
  INV_X1 U560 ( .A(initial_mask_in[31]), .ZN(n368) );
  OAI22_X1 U561 ( .A1(n81), .A2(n852), .B1(n90), .B2(n369), .ZN(n1044) );
  INV_X1 U562 ( .A(next_pc_in[0]), .ZN(n369) );
  OAI22_X1 U563 ( .A1(n81), .A2(n851), .B1(n90), .B2(n370), .ZN(n1043) );
  INV_X1 U564 ( .A(next_pc_in[1]), .ZN(n370) );
  OAI22_X1 U565 ( .A1(n81), .A2(n850), .B1(n90), .B2(n371), .ZN(n1042) );
  INV_X1 U566 ( .A(next_pc_in[2]), .ZN(n371) );
  OAI22_X1 U567 ( .A1(n81), .A2(n849), .B1(n90), .B2(n372), .ZN(n1041) );
  INV_X1 U568 ( .A(next_pc_in[3]), .ZN(n372) );
  OAI22_X1 U569 ( .A1(n81), .A2(n848), .B1(n90), .B2(n373), .ZN(n1040) );
  INV_X1 U570 ( .A(next_pc_in[4]), .ZN(n373) );
  OAI22_X1 U571 ( .A1(n81), .A2(n847), .B1(n90), .B2(n374), .ZN(n1039) );
  INV_X1 U572 ( .A(next_pc_in[5]), .ZN(n374) );
  OAI22_X1 U573 ( .A1(n81), .A2(n846), .B1(n90), .B2(n375), .ZN(n1038) );
  INV_X1 U574 ( .A(next_pc_in[6]), .ZN(n375) );
  OAI22_X1 U575 ( .A1(n81), .A2(n845), .B1(n90), .B2(n376), .ZN(n1037) );
  INV_X1 U576 ( .A(next_pc_in[7]), .ZN(n376) );
  OAI22_X1 U577 ( .A1(n81), .A2(n844), .B1(n90), .B2(n377), .ZN(n1036) );
  INV_X1 U578 ( .A(next_pc_in[8]), .ZN(n377) );
  OAI22_X1 U579 ( .A1(n81), .A2(n843), .B1(n90), .B2(n378), .ZN(n1035) );
  INV_X1 U580 ( .A(next_pc_in[9]), .ZN(n378) );
  OAI22_X1 U581 ( .A1(n81), .A2(n842), .B1(n91), .B2(n379), .ZN(n1034) );
  INV_X1 U582 ( .A(next_pc_in[10]), .ZN(n379) );
  OAI22_X1 U583 ( .A1(n81), .A2(n841), .B1(n91), .B2(n380), .ZN(n1033) );
  INV_X1 U584 ( .A(next_pc_in[11]), .ZN(n380) );
  OAI22_X1 U585 ( .A1(n80), .A2(n840), .B1(n91), .B2(n381), .ZN(n1032) );
  INV_X1 U586 ( .A(next_pc_in[12]), .ZN(n381) );
  OAI22_X1 U587 ( .A1(n77), .A2(n839), .B1(n91), .B2(n382), .ZN(n1031) );
  INV_X1 U588 ( .A(next_pc_in[13]), .ZN(n382) );
  OAI22_X1 U589 ( .A1(n79), .A2(n838), .B1(n91), .B2(n383), .ZN(n1030) );
  INV_X1 U590 ( .A(next_pc_in[14]), .ZN(n383) );
  OAI22_X1 U591 ( .A1(n82), .A2(n837), .B1(n91), .B2(n384), .ZN(n1029) );
  INV_X1 U592 ( .A(next_pc_in[15]), .ZN(n384) );
  OAI22_X1 U593 ( .A1(n81), .A2(n836), .B1(n91), .B2(n385), .ZN(n1028) );
  INV_X1 U594 ( .A(next_pc_in[16]), .ZN(n385) );
  OAI22_X1 U595 ( .A1(n80), .A2(n835), .B1(n91), .B2(n386), .ZN(n1027) );
  INV_X1 U596 ( .A(next_pc_in[17]), .ZN(n386) );
  OAI22_X1 U597 ( .A1(n77), .A2(n834), .B1(n91), .B2(n387), .ZN(n1026) );
  INV_X1 U598 ( .A(next_pc_in[18]), .ZN(n387) );
  OAI22_X1 U599 ( .A1(n79), .A2(n833), .B1(n91), .B2(n388), .ZN(n1025) );
  INV_X1 U600 ( .A(next_pc_in[19]), .ZN(n388) );
  OAI22_X1 U601 ( .A1(n82), .A2(n832), .B1(n91), .B2(n389), .ZN(n1024) );
  INV_X1 U602 ( .A(next_pc_in[20]), .ZN(n389) );
  OAI22_X1 U603 ( .A1(n81), .A2(n831), .B1(n91), .B2(n390), .ZN(n1023) );
  INV_X1 U604 ( .A(next_pc_in[21]), .ZN(n390) );
  OAI22_X1 U605 ( .A1(n80), .A2(n830), .B1(n92), .B2(n391), .ZN(n1022) );
  INV_X1 U606 ( .A(next_pc_in[22]), .ZN(n391) );
  OAI22_X1 U607 ( .A1(n82), .A2(n829), .B1(n92), .B2(n392), .ZN(n1021) );
  INV_X1 U608 ( .A(next_pc_in[23]), .ZN(n392) );
  OAI22_X1 U609 ( .A1(n82), .A2(n828), .B1(n92), .B2(n393), .ZN(n1020) );
  INV_X1 U610 ( .A(next_pc_in[24]), .ZN(n393) );
  OAI22_X1 U611 ( .A1(n82), .A2(n827), .B1(n92), .B2(n394), .ZN(n1019) );
  INV_X1 U612 ( .A(next_pc_in[25]), .ZN(n394) );
  OAI22_X1 U613 ( .A1(n82), .A2(n826), .B1(n92), .B2(n395), .ZN(n1018) );
  INV_X1 U614 ( .A(next_pc_in[26]), .ZN(n395) );
  OAI22_X1 U615 ( .A1(n82), .A2(n825), .B1(n92), .B2(n396), .ZN(n1017) );
  INV_X1 U616 ( .A(next_pc_in[27]), .ZN(n396) );
  OAI22_X1 U617 ( .A1(n82), .A2(n824), .B1(n92), .B2(n397), .ZN(n1016) );
  INV_X1 U618 ( .A(next_pc_in[28]), .ZN(n397) );
  OAI22_X1 U619 ( .A1(n82), .A2(n823), .B1(n92), .B2(n398), .ZN(n1015) );
  INV_X1 U620 ( .A(next_pc_in[29]), .ZN(n398) );
  OAI22_X1 U621 ( .A1(n82), .A2(n822), .B1(n92), .B2(n399), .ZN(n1014) );
  INV_X1 U622 ( .A(next_pc_in[30]), .ZN(n399) );
  OAI22_X1 U623 ( .A1(n82), .A2(n821), .B1(n92), .B2(n400), .ZN(n1013) );
  INV_X1 U624 ( .A(next_pc_in[31]), .ZN(n400) );
  OAI22_X1 U625 ( .A1(n82), .A2(n820), .B1(n92), .B2(n401), .ZN(n1012) );
  INV_X1 U626 ( .A(gprs_base_addr_in[0]), .ZN(n401) );
  OAI22_X1 U627 ( .A1(n82), .A2(n819), .B1(n92), .B2(n402), .ZN(n1011) );
  INV_X1 U628 ( .A(gprs_base_addr_in[1]), .ZN(n402) );
  OAI22_X1 U629 ( .A1(n81), .A2(n818), .B1(n93), .B2(n403), .ZN(n1010) );
  INV_X1 U630 ( .A(gprs_base_addr_in[2]), .ZN(n403) );
  OAI22_X1 U631 ( .A1(n82), .A2(n817), .B1(n93), .B2(n404), .ZN(n1009) );
  INV_X1 U632 ( .A(gprs_base_addr_in[3]), .ZN(n404) );
  OAI22_X1 U633 ( .A1(n82), .A2(n816), .B1(n93), .B2(n405), .ZN(n1008) );
  INV_X1 U634 ( .A(gprs_base_addr_in[4]), .ZN(n405) );
  OAI22_X1 U635 ( .A1(n80), .A2(n815), .B1(n93), .B2(n406), .ZN(n1007) );
  INV_X1 U636 ( .A(gprs_base_addr_in[5]), .ZN(n406) );
  OAI22_X1 U637 ( .A1(n78), .A2(n814), .B1(n93), .B2(n407), .ZN(n1006) );
  INV_X1 U638 ( .A(gprs_base_addr_in[6]), .ZN(n407) );
  OAI22_X1 U639 ( .A1(n82), .A2(n813), .B1(n93), .B2(n408), .ZN(n1005) );
  INV_X1 U640 ( .A(gprs_base_addr_in[7]), .ZN(n408) );
  OAI22_X1 U641 ( .A1(n79), .A2(n812), .B1(n93), .B2(n409), .ZN(n1004) );
  INV_X1 U642 ( .A(gprs_base_addr_in[8]), .ZN(n409) );
  OAI22_X1 U643 ( .A1(n77), .A2(n811), .B1(n93), .B2(n410), .ZN(n1003) );
  INV_X1 U644 ( .A(shmem_base_addr_in[0]), .ZN(n410) );
  OAI22_X1 U645 ( .A1(n78), .A2(n810), .B1(n93), .B2(n411), .ZN(n1002) );
  INV_X1 U646 ( .A(shmem_base_addr_in[1]), .ZN(n411) );
  OAI22_X1 U647 ( .A1(n77), .A2(n809), .B1(n93), .B2(n412), .ZN(n1001) );
  INV_X1 U648 ( .A(shmem_base_addr_in[2]), .ZN(n412) );
  OAI22_X1 U649 ( .A1(n77), .A2(n808), .B1(n83), .B2(n413), .ZN(n1000) );
  INV_X1 U650 ( .A(shmem_base_addr_in[3]), .ZN(n413) );
  NAND2_X1 U651 ( .A1(n181), .A2(n78), .ZN(n149) );
  NOR2_X1 U652 ( .A1(n304), .A2(n102), .ZN(n181) );
  OAI21_X1 U653 ( .B1(n182), .B2(n304), .A(n99), .ZN(n414) );
  INV_X1 U654 ( .A(en), .ZN(n304) );
  INV_X1 U655 ( .A(n302), .ZN(n182) );
  NAND2_X1 U656 ( .A1(warp_lane_id_in[1]), .A2(warp_lane_id_in[0]), .ZN(n302)
         );
  INV_X1 U657 ( .A(n257), .ZN(n187) );
  NOR3_X1 U658 ( .A1(warp_checker_state_machine[1]), .A2(
        warp_checker_state_machine[2]), .A3(n3), .ZN(n257) );
  INV_X1 U659 ( .A(n190), .ZN(n197) );
  NOR3_X1 U660 ( .A1(warp_checker_state_machine[0]), .A2(
        warp_checker_state_machine[1]), .A3(n8), .ZN(n190) );
  NOR2_X1 U661 ( .A1(n415), .A2(n416), .ZN(fence_id_mask[9]) );
  INV_X1 U662 ( .A(fence_regs_fence_en_in[9]), .ZN(n415) );
  NOR2_X1 U663 ( .A1(n417), .A2(n418), .ZN(fence_id_mask[8]) );
  INV_X1 U664 ( .A(fence_regs_fence_en_in[8]), .ZN(n417) );
  NOR2_X1 U665 ( .A1(n419), .A2(n420), .ZN(fence_id_mask[7]) );
  INV_X1 U666 ( .A(fence_regs_fence_en_in[7]), .ZN(n419) );
  NOR2_X1 U667 ( .A1(n421), .A2(n422), .ZN(fence_id_mask[6]) );
  INV_X1 U668 ( .A(fence_regs_fence_en_in[6]), .ZN(n421) );
  NOR2_X1 U669 ( .A1(n423), .A2(n424), .ZN(fence_id_mask[5]) );
  INV_X1 U670 ( .A(fence_regs_fence_en_in[5]), .ZN(n423) );
  NOR2_X1 U671 ( .A1(n425), .A2(n426), .ZN(fence_id_mask[4]) );
  INV_X1 U672 ( .A(fence_regs_fence_en_in[4]), .ZN(n425) );
  NOR2_X1 U673 ( .A1(n427), .A2(n428), .ZN(fence_id_mask[3]) );
  INV_X1 U674 ( .A(fence_regs_fence_en_in[3]), .ZN(n427) );
  NOR2_X1 U675 ( .A1(n429), .A2(n430), .ZN(fence_id_mask[31]) );
  INV_X1 U676 ( .A(fence_regs_fence_en_in[31]), .ZN(n429) );
  NOR2_X1 U677 ( .A1(n431), .A2(n432), .ZN(fence_id_mask[30]) );
  INV_X1 U678 ( .A(fence_regs_fence_en_in[30]), .ZN(n431) );
  NOR2_X1 U679 ( .A1(n433), .A2(n434), .ZN(fence_id_mask[2]) );
  INV_X1 U680 ( .A(fence_regs_fence_en_in[2]), .ZN(n433) );
  NOR2_X1 U681 ( .A1(n435), .A2(n436), .ZN(fence_id_mask[29]) );
  INV_X1 U682 ( .A(fence_regs_fence_en_in[29]), .ZN(n435) );
  NOR2_X1 U683 ( .A1(n437), .A2(n438), .ZN(fence_id_mask[28]) );
  INV_X1 U684 ( .A(fence_regs_fence_en_in[28]), .ZN(n437) );
  NOR2_X1 U685 ( .A1(n439), .A2(n440), .ZN(fence_id_mask[27]) );
  INV_X1 U686 ( .A(fence_regs_fence_en_in[27]), .ZN(n439) );
  NOR2_X1 U687 ( .A1(n441), .A2(n442), .ZN(fence_id_mask[26]) );
  INV_X1 U688 ( .A(fence_regs_fence_en_in[26]), .ZN(n441) );
  NOR2_X1 U689 ( .A1(n443), .A2(n444), .ZN(fence_id_mask[25]) );
  INV_X1 U690 ( .A(fence_regs_fence_en_in[25]), .ZN(n443) );
  NOR2_X1 U691 ( .A1(n445), .A2(n446), .ZN(fence_id_mask[24]) );
  INV_X1 U692 ( .A(fence_regs_fence_en_in[24]), .ZN(n445) );
  NOR2_X1 U693 ( .A1(n447), .A2(n448), .ZN(fence_id_mask[23]) );
  INV_X1 U694 ( .A(fence_regs_fence_en_in[23]), .ZN(n447) );
  NOR2_X1 U695 ( .A1(n449), .A2(n450), .ZN(fence_id_mask[22]) );
  INV_X1 U696 ( .A(fence_regs_fence_en_in[22]), .ZN(n449) );
  NOR2_X1 U697 ( .A1(n451), .A2(n452), .ZN(fence_id_mask[21]) );
  INV_X1 U698 ( .A(fence_regs_fence_en_in[21]), .ZN(n451) );
  NOR2_X1 U699 ( .A1(n453), .A2(n454), .ZN(fence_id_mask[20]) );
  INV_X1 U700 ( .A(fence_regs_fence_en_in[20]), .ZN(n453) );
  NOR2_X1 U701 ( .A1(n455), .A2(n456), .ZN(fence_id_mask[1]) );
  INV_X1 U702 ( .A(fence_regs_fence_en_in[1]), .ZN(n455) );
  NOR2_X1 U703 ( .A1(n457), .A2(n458), .ZN(fence_id_mask[19]) );
  INV_X1 U704 ( .A(fence_regs_fence_en_in[19]), .ZN(n457) );
  NOR2_X1 U705 ( .A1(n459), .A2(n460), .ZN(fence_id_mask[18]) );
  INV_X1 U706 ( .A(fence_regs_fence_en_in[18]), .ZN(n459) );
  NOR2_X1 U707 ( .A1(n461), .A2(n462), .ZN(fence_id_mask[17]) );
  INV_X1 U708 ( .A(fence_regs_fence_en_in[17]), .ZN(n461) );
  NOR2_X1 U709 ( .A1(n463), .A2(n464), .ZN(fence_id_mask[16]) );
  INV_X1 U710 ( .A(fence_regs_fence_en_in[16]), .ZN(n463) );
  NOR2_X1 U711 ( .A1(n465), .A2(n466), .ZN(fence_id_mask[15]) );
  INV_X1 U712 ( .A(fence_regs_fence_en_in[15]), .ZN(n465) );
  NOR2_X1 U713 ( .A1(n467), .A2(n468), .ZN(fence_id_mask[14]) );
  INV_X1 U714 ( .A(fence_regs_fence_en_in[14]), .ZN(n467) );
  NOR2_X1 U715 ( .A1(n469), .A2(n470), .ZN(fence_id_mask[13]) );
  INV_X1 U716 ( .A(fence_regs_fence_en_in[13]), .ZN(n469) );
  NOR2_X1 U717 ( .A1(n471), .A2(n472), .ZN(fence_id_mask[12]) );
  INV_X1 U718 ( .A(fence_regs_fence_en_in[12]), .ZN(n471) );
  NOR2_X1 U719 ( .A1(n473), .A2(n474), .ZN(fence_id_mask[11]) );
  INV_X1 U720 ( .A(fence_regs_fence_en_in[11]), .ZN(n473) );
  NOR2_X1 U721 ( .A1(n475), .A2(n476), .ZN(fence_id_mask[10]) );
  INV_X1 U722 ( .A(fence_regs_fence_en_in[10]), .ZN(n475) );
  NOR2_X1 U723 ( .A1(n477), .A2(n478), .ZN(fence_id_mask[0]) );
  INV_X1 U724 ( .A(fence_regs_fence_en_in[0]), .ZN(n477) );
  AOI21_X1 U725 ( .B1(n479), .B2(n480), .A(n416), .ZN(cta_id_mask_rev[9]) );
  NAND4_X1 U726 ( .A1(n481), .A2(n482), .A3(n483), .A4(n484), .ZN(n416) );
  XNOR2_X1 U727 ( .A(n137), .B(\fence_regs_cta_id_in[9><0] ), .ZN(n484) );
  XNOR2_X1 U728 ( .A(n139), .B(\fence_regs_cta_id_in[9><1] ), .ZN(n483) );
  XNOR2_X1 U729 ( .A(n141), .B(\fence_regs_cta_id_in[9><2] ), .ZN(n482) );
  XNOR2_X1 U730 ( .A(n143), .B(\fence_regs_cta_id_in[9><3] ), .ZN(n481) );
  AOI21_X1 U731 ( .B1(n479), .B2(n485), .A(n418), .ZN(cta_id_mask_rev[8]) );
  NAND4_X1 U732 ( .A1(n486), .A2(n487), .A3(n488), .A4(n489), .ZN(n418) );
  XNOR2_X1 U733 ( .A(n137), .B(\fence_regs_cta_id_in[8><0] ), .ZN(n489) );
  XNOR2_X1 U734 ( .A(n139), .B(\fence_regs_cta_id_in[8><1] ), .ZN(n488) );
  XNOR2_X1 U735 ( .A(n141), .B(\fence_regs_cta_id_in[8><2] ), .ZN(n487) );
  XNOR2_X1 U736 ( .A(n143), .B(\fence_regs_cta_id_in[8><3] ), .ZN(n486) );
  NOR2_X1 U737 ( .A1(n490), .A2(n420), .ZN(cta_id_mask_rev[7]) );
  NAND4_X1 U738 ( .A1(n491), .A2(n492), .A3(n493), .A4(n494), .ZN(n420) );
  XNOR2_X1 U739 ( .A(n137), .B(\fence_regs_cta_id_in[7><0] ), .ZN(n494) );
  XNOR2_X1 U740 ( .A(n139), .B(\fence_regs_cta_id_in[7><1] ), .ZN(n493) );
  XNOR2_X1 U741 ( .A(n141), .B(\fence_regs_cta_id_in[7><2] ), .ZN(n492) );
  XNOR2_X1 U742 ( .A(n143), .B(\fence_regs_cta_id_in[7><3] ), .ZN(n491) );
  NOR2_X1 U743 ( .A1(n495), .A2(n422), .ZN(cta_id_mask_rev[6]) );
  NAND4_X1 U744 ( .A1(n496), .A2(n497), .A3(n498), .A4(n499), .ZN(n422) );
  XNOR2_X1 U745 ( .A(n137), .B(\fence_regs_cta_id_in[6><0] ), .ZN(n499) );
  XNOR2_X1 U746 ( .A(n139), .B(\fence_regs_cta_id_in[6><1] ), .ZN(n498) );
  XNOR2_X1 U747 ( .A(n141), .B(\fence_regs_cta_id_in[6><2] ), .ZN(n497) );
  XNOR2_X1 U748 ( .A(n143), .B(\fence_regs_cta_id_in[6><3] ), .ZN(n496) );
  AOI21_X1 U749 ( .B1(n500), .B2(warps_per_block_in[2]), .A(n501), .ZN(n495)
         );
  NOR2_X1 U750 ( .A1(n502), .A2(n424), .ZN(cta_id_mask_rev[5]) );
  NAND4_X1 U751 ( .A1(n503), .A2(n504), .A3(n505), .A4(n506), .ZN(n424) );
  XNOR2_X1 U752 ( .A(n137), .B(\fence_regs_cta_id_in[5><0] ), .ZN(n506) );
  XNOR2_X1 U753 ( .A(n139), .B(\fence_regs_cta_id_in[5><1] ), .ZN(n505) );
  XNOR2_X1 U754 ( .A(n141), .B(\fence_regs_cta_id_in[5><2] ), .ZN(n504) );
  XNOR2_X1 U755 ( .A(n143), .B(\fence_regs_cta_id_in[5><3] ), .ZN(n503) );
  AOI21_X1 U756 ( .B1(warps_per_block_in[2]), .B2(warps_per_block_in[1]), .A(
        n501), .ZN(n502) );
  NOR2_X1 U757 ( .A1(n507), .A2(n426), .ZN(cta_id_mask_rev[4]) );
  NAND4_X1 U758 ( .A1(n508), .A2(n509), .A3(n510), .A4(n511), .ZN(n426) );
  XNOR2_X1 U759 ( .A(n137), .B(\fence_regs_cta_id_in[4><0] ), .ZN(n511) );
  XNOR2_X1 U760 ( .A(n139), .B(\fence_regs_cta_id_in[4><1] ), .ZN(n510) );
  XNOR2_X1 U761 ( .A(n141), .B(\fence_regs_cta_id_in[4><2] ), .ZN(n509) );
  XNOR2_X1 U762 ( .A(n143), .B(\fence_regs_cta_id_in[4><3] ), .ZN(n508) );
  AOI21_X1 U763 ( .B1(warps_per_block_in[2]), .B2(n512), .A(n501), .ZN(n507)
         );
  NOR2_X1 U764 ( .A1(n513), .A2(n428), .ZN(cta_id_mask_rev[3]) );
  NAND4_X1 U765 ( .A1(n514), .A2(n515), .A3(n516), .A4(n517), .ZN(n428) );
  XNOR2_X1 U766 ( .A(n137), .B(\fence_regs_cta_id_in[3><0] ), .ZN(n517) );
  XNOR2_X1 U767 ( .A(n139), .B(\fence_regs_cta_id_in[3><1] ), .ZN(n516) );
  XNOR2_X1 U768 ( .A(n141), .B(\fence_regs_cta_id_in[3><2] ), .ZN(n515) );
  XNOR2_X1 U769 ( .A(n143), .B(\fence_regs_cta_id_in[3><3] ), .ZN(n514) );
  NOR2_X1 U770 ( .A1(n518), .A2(n430), .ZN(cta_id_mask_rev[31]) );
  NAND4_X1 U771 ( .A1(n519), .A2(n520), .A3(n521), .A4(n522), .ZN(n430) );
  XNOR2_X1 U772 ( .A(n137), .B(\fence_regs_cta_id_in[31><0] ), .ZN(n522) );
  XNOR2_X1 U773 ( .A(n139), .B(\fence_regs_cta_id_in[31><1] ), .ZN(n521) );
  XNOR2_X1 U774 ( .A(n141), .B(\fence_regs_cta_id_in[31><2] ), .ZN(n520) );
  XNOR2_X1 U775 ( .A(n143), .B(\fence_regs_cta_id_in[31><3] ), .ZN(n519) );
  AOI21_X1 U776 ( .B1(n518), .B2(n523), .A(n432), .ZN(cta_id_mask_rev[30]) );
  NAND4_X1 U777 ( .A1(n524), .A2(n525), .A3(n526), .A4(n527), .ZN(n432) );
  XNOR2_X1 U778 ( .A(n137), .B(\fence_regs_cta_id_in[30><0] ), .ZN(n527) );
  XNOR2_X1 U779 ( .A(n139), .B(\fence_regs_cta_id_in[30><1] ), .ZN(n526) );
  XNOR2_X1 U780 ( .A(n141), .B(\fence_regs_cta_id_in[30><2] ), .ZN(n525) );
  XNOR2_X1 U781 ( .A(n143), .B(\fence_regs_cta_id_in[30><3] ), .ZN(n524) );
  NAND3_X1 U782 ( .A1(n528), .A2(warps_per_block_in[0]), .A3(n529), .ZN(n523)
         );
  AOI21_X1 U783 ( .B1(n530), .B2(n490), .A(n434), .ZN(cta_id_mask_rev[2]) );
  NAND4_X1 U784 ( .A1(n531), .A2(n532), .A3(n533), .A4(n534), .ZN(n434) );
  XNOR2_X1 U785 ( .A(n137), .B(\fence_regs_cta_id_in[2><0] ), .ZN(n534) );
  XNOR2_X1 U786 ( .A(n139), .B(\fence_regs_cta_id_in[2><1] ), .ZN(n533) );
  XNOR2_X1 U787 ( .A(n141), .B(\fence_regs_cta_id_in[2><2] ), .ZN(n532) );
  XNOR2_X1 U788 ( .A(n143), .B(\fence_regs_cta_id_in[2><3] ), .ZN(n531) );
  NOR2_X1 U789 ( .A1(n535), .A2(n436), .ZN(cta_id_mask_rev[29]) );
  NAND4_X1 U790 ( .A1(n536), .A2(n537), .A3(n538), .A4(n539), .ZN(n436) );
  XNOR2_X1 U791 ( .A(n137), .B(\fence_regs_cta_id_in[29><0] ), .ZN(n539) );
  XNOR2_X1 U792 ( .A(n139), .B(\fence_regs_cta_id_in[29><1] ), .ZN(n538) );
  XNOR2_X1 U793 ( .A(n141), .B(\fence_regs_cta_id_in[29><2] ), .ZN(n537) );
  XNOR2_X1 U794 ( .A(n143), .B(\fence_regs_cta_id_in[29><3] ), .ZN(n536) );
  AOI21_X1 U795 ( .B1(n529), .B2(n528), .A(n540), .ZN(n535) );
  NOR2_X1 U796 ( .A1(n541), .A2(n438), .ZN(cta_id_mask_rev[28]) );
  NAND4_X1 U797 ( .A1(n542), .A2(n543), .A3(n544), .A4(n545), .ZN(n438) );
  XNOR2_X1 U798 ( .A(n137), .B(\fence_regs_cta_id_in[28><0] ), .ZN(n545) );
  XNOR2_X1 U799 ( .A(n139), .B(\fence_regs_cta_id_in[28><1] ), .ZN(n544) );
  XNOR2_X1 U800 ( .A(n141), .B(\fence_regs_cta_id_in[28><2] ), .ZN(n543) );
  XNOR2_X1 U801 ( .A(n143), .B(\fence_regs_cta_id_in[28><3] ), .ZN(n542) );
  AOI21_X1 U802 ( .B1(n546), .B2(n529), .A(n540), .ZN(n541) );
  NOR2_X1 U803 ( .A1(n547), .A2(n440), .ZN(cta_id_mask_rev[27]) );
  NAND4_X1 U804 ( .A1(n548), .A2(n549), .A3(n550), .A4(n551), .ZN(n440) );
  XNOR2_X1 U805 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[27><0] ), .ZN(
        n551) );
  XNOR2_X1 U806 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[27><1] ), .ZN(
        n550) );
  XNOR2_X1 U807 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[27><2] ), .ZN(
        n549) );
  XNOR2_X1 U808 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[27><3] ), .ZN(
        n548) );
  AOI21_X1 U809 ( .B1(n518), .B2(n552), .A(n442), .ZN(cta_id_mask_rev[26]) );
  NAND4_X1 U810 ( .A1(n553), .A2(n554), .A3(n555), .A4(n556), .ZN(n442) );
  XNOR2_X1 U811 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[26><0] ), .ZN(
        n556) );
  XNOR2_X1 U812 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[26><1] ), .ZN(
        n555) );
  XNOR2_X1 U813 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[26><2] ), .ZN(
        n554) );
  XNOR2_X1 U814 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[26><3] ), .ZN(
        n553) );
  NAND3_X1 U815 ( .A1(warps_per_block_in[3]), .A2(n557), .A3(
        warps_per_block_in[4]), .ZN(n552) );
  INV_X1 U816 ( .A(n540), .ZN(n518) );
  AOI21_X1 U817 ( .B1(n547), .B2(n558), .A(n444), .ZN(cta_id_mask_rev[25]) );
  NAND4_X1 U818 ( .A1(n559), .A2(n560), .A3(n561), .A4(n562), .ZN(n444) );
  XNOR2_X1 U819 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[25><0] ), .ZN(
        n562) );
  XNOR2_X1 U820 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[25><1] ), .ZN(
        n561) );
  XNOR2_X1 U821 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[25><2] ), .ZN(
        n560) );
  XNOR2_X1 U822 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[25><3] ), .ZN(
        n559) );
  NAND2_X1 U823 ( .A1(n528), .A2(warps_per_block_in[4]), .ZN(n558) );
  AOI21_X1 U824 ( .B1(n547), .B2(n563), .A(n446), .ZN(cta_id_mask_rev[24]) );
  NAND4_X1 U825 ( .A1(n564), .A2(n565), .A3(n566), .A4(n567), .ZN(n446) );
  XNOR2_X1 U826 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[24><0] ), .ZN(
        n567) );
  XNOR2_X1 U827 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[24><1] ), .ZN(
        n566) );
  XNOR2_X1 U828 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[24><2] ), .ZN(
        n565) );
  XNOR2_X1 U829 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[24><3] ), .ZN(
        n564) );
  NAND2_X1 U830 ( .A1(n546), .A2(warps_per_block_in[4]), .ZN(n563) );
  AOI21_X1 U831 ( .B1(warps_per_block_in[3]), .B2(n529), .A(n540), .ZN(n547)
         );
  NOR2_X1 U832 ( .A1(n568), .A2(n448), .ZN(cta_id_mask_rev[23]) );
  NAND4_X1 U833 ( .A1(n569), .A2(n570), .A3(n571), .A4(n572), .ZN(n448) );
  XNOR2_X1 U834 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[23><0] ), .ZN(
        n572) );
  XNOR2_X1 U835 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[23><1] ), .ZN(
        n571) );
  XNOR2_X1 U836 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[23><2] ), .ZN(
        n570) );
  XNOR2_X1 U837 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[23><3] ), .ZN(
        n569) );
  AOI21_X1 U838 ( .B1(n568), .B2(n573), .A(n450), .ZN(cta_id_mask_rev[22]) );
  NAND4_X1 U839 ( .A1(n574), .A2(n575), .A3(n576), .A4(n577), .ZN(n450) );
  XNOR2_X1 U840 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[22><0] ), .ZN(
        n577) );
  XNOR2_X1 U841 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[22><1] ), .ZN(
        n576) );
  XNOR2_X1 U842 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[22><2] ), .ZN(
        n575) );
  XNOR2_X1 U843 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[22><3] ), .ZN(
        n574) );
  NAND2_X1 U844 ( .A1(n529), .A2(n500), .ZN(n573) );
  AOI21_X1 U845 ( .B1(n568), .B2(n578), .A(n452), .ZN(cta_id_mask_rev[21]) );
  NAND4_X1 U846 ( .A1(n579), .A2(n580), .A3(n581), .A4(n582), .ZN(n452) );
  XNOR2_X1 U847 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[21><0] ), .ZN(
        n582) );
  XNOR2_X1 U848 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[21><1] ), .ZN(
        n581) );
  XNOR2_X1 U849 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[21><2] ), .ZN(
        n580) );
  XNOR2_X1 U850 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[21><3] ), .ZN(
        n579) );
  NAND2_X1 U851 ( .A1(n529), .A2(warps_per_block_in[1]), .ZN(n578) );
  AOI21_X1 U852 ( .B1(n568), .B2(n583), .A(n454), .ZN(cta_id_mask_rev[20]) );
  NAND4_X1 U853 ( .A1(n584), .A2(n585), .A3(n586), .A4(n587), .ZN(n454) );
  XNOR2_X1 U854 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[20><0] ), .ZN(
        n587) );
  XNOR2_X1 U855 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[20><1] ), .ZN(
        n586) );
  XNOR2_X1 U856 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[20><2] ), .ZN(
        n585) );
  XNOR2_X1 U857 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[20><3] ), .ZN(
        n584) );
  NAND2_X1 U858 ( .A1(n529), .A2(n512), .ZN(n583) );
  INV_X1 U859 ( .A(n588), .ZN(n529) );
  AOI21_X1 U860 ( .B1(n513), .B2(n589), .A(n456), .ZN(cta_id_mask_rev[1]) );
  NAND4_X1 U861 ( .A1(n590), .A2(n591), .A3(n592), .A4(n593), .ZN(n456) );
  XNOR2_X1 U862 ( .A(n137), .B(\fence_regs_cta_id_in[1><0] ), .ZN(n593) );
  XNOR2_X1 U863 ( .A(n139), .B(\fence_regs_cta_id_in[1><1] ), .ZN(n592) );
  XNOR2_X1 U864 ( .A(n141), .B(\fence_regs_cta_id_in[1><2] ), .ZN(n591) );
  XNOR2_X1 U865 ( .A(n143), .B(\fence_regs_cta_id_in[1><3] ), .ZN(n590) );
  INV_X1 U866 ( .A(warps_per_block_in[1]), .ZN(n589) );
  NOR2_X1 U867 ( .A1(n594), .A2(n458), .ZN(cta_id_mask_rev[19]) );
  NAND4_X1 U868 ( .A1(n595), .A2(n596), .A3(n597), .A4(n598), .ZN(n458) );
  XNOR2_X1 U869 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[19><0] ), .ZN(
        n598) );
  XNOR2_X1 U870 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[19><1] ), .ZN(
        n597) );
  XNOR2_X1 U871 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[19><2] ), .ZN(
        n596) );
  XNOR2_X1 U872 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[19><3] ), .ZN(
        n595) );
  INV_X1 U873 ( .A(n599), .ZN(n594) );
  AOI21_X1 U874 ( .B1(n568), .B2(n600), .A(n460), .ZN(cta_id_mask_rev[18]) );
  NAND4_X1 U875 ( .A1(n601), .A2(n602), .A3(n603), .A4(n604), .ZN(n460) );
  XNOR2_X1 U876 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[18><0] ), .ZN(
        n604) );
  XNOR2_X1 U877 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[18><1] ), .ZN(
        n603) );
  XNOR2_X1 U878 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[18><2] ), .ZN(
        n602) );
  XNOR2_X1 U879 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[18><3] ), .ZN(
        n601) );
  NAND2_X1 U880 ( .A1(warps_per_block_in[4]), .A2(n557), .ZN(n600) );
  NOR2_X1 U881 ( .A1(n605), .A2(n462), .ZN(cta_id_mask_rev[17]) );
  NAND4_X1 U882 ( .A1(n606), .A2(n607), .A3(n608), .A4(n609), .ZN(n462) );
  XNOR2_X1 U883 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[17><0] ), .ZN(
        n609) );
  XNOR2_X1 U884 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[17><1] ), .ZN(
        n608) );
  XNOR2_X1 U885 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[17><2] ), .ZN(
        n607) );
  XNOR2_X1 U886 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[17><3] ), .ZN(
        n606) );
  AOI21_X1 U887 ( .B1(warps_per_block_in[4]), .B2(warps_per_block_in[1]), .A(
        n599), .ZN(n605) );
  NOR2_X1 U888 ( .A1(n610), .A2(n464), .ZN(cta_id_mask_rev[16]) );
  NAND4_X1 U889 ( .A1(n611), .A2(n612), .A3(n613), .A4(n614), .ZN(n464) );
  XNOR2_X1 U890 ( .A(n137), .B(\fence_regs_cta_id_in[16><0] ), .ZN(n614) );
  XNOR2_X1 U891 ( .A(n139), .B(\fence_regs_cta_id_in[16><1] ), .ZN(n613) );
  XNOR2_X1 U892 ( .A(n141), .B(\fence_regs_cta_id_in[16><2] ), .ZN(n612) );
  XNOR2_X1 U893 ( .A(n143), .B(\fence_regs_cta_id_in[16><3] ), .ZN(n611) );
  AOI21_X1 U894 ( .B1(warps_per_block_in[4]), .B2(n512), .A(n599), .ZN(n610)
         );
  NAND2_X1 U895 ( .A1(n568), .A2(n588), .ZN(n599) );
  NAND2_X1 U896 ( .A1(warps_per_block_in[4]), .A2(warps_per_block_in[2]), .ZN(
        n588) );
  AOI21_X1 U897 ( .B1(warps_per_block_in[3]), .B2(warps_per_block_in[4]), .A(
        n540), .ZN(n568) );
  NOR2_X1 U898 ( .A1(n615), .A2(n466), .ZN(cta_id_mask_rev[15]) );
  NAND4_X1 U899 ( .A1(n616), .A2(n617), .A3(n618), .A4(n619), .ZN(n466) );
  XNOR2_X1 U900 ( .A(n137), .B(\fence_regs_cta_id_in[15><0] ), .ZN(n619) );
  XNOR2_X1 U901 ( .A(n139), .B(\fence_regs_cta_id_in[15><1] ), .ZN(n618) );
  XNOR2_X1 U902 ( .A(n141), .B(\fence_regs_cta_id_in[15><2] ), .ZN(n617) );
  XNOR2_X1 U903 ( .A(n143), .B(\fence_regs_cta_id_in[15><3] ), .ZN(n616) );
  AOI21_X1 U904 ( .B1(n615), .B2(n620), .A(n468), .ZN(cta_id_mask_rev[14]) );
  NAND4_X1 U905 ( .A1(n621), .A2(n622), .A3(n623), .A4(n624), .ZN(n468) );
  XNOR2_X1 U906 ( .A(n137), .B(\fence_regs_cta_id_in[14><0] ), .ZN(n624) );
  XNOR2_X1 U907 ( .A(n139), .B(\fence_regs_cta_id_in[14><1] ), .ZN(n623) );
  XNOR2_X1 U908 ( .A(n141), .B(\fence_regs_cta_id_in[14><2] ), .ZN(n622) );
  XNOR2_X1 U909 ( .A(n143), .B(\fence_regs_cta_id_in[14><3] ), .ZN(n621) );
  NAND3_X1 U910 ( .A1(warps_per_block_in[0]), .A2(warps_per_block_in[2]), .A3(
        n528), .ZN(n620) );
  AOI21_X1 U911 ( .B1(n615), .B2(n625), .A(n470), .ZN(cta_id_mask_rev[13]) );
  NAND4_X1 U912 ( .A1(n626), .A2(n627), .A3(n628), .A4(n629), .ZN(n470) );
  XNOR2_X1 U913 ( .A(n137), .B(\fence_regs_cta_id_in[13><0] ), .ZN(n629) );
  XNOR2_X1 U914 ( .A(n139), .B(\fence_regs_cta_id_in[13><1] ), .ZN(n628) );
  XNOR2_X1 U915 ( .A(n141), .B(\fence_regs_cta_id_in[13><2] ), .ZN(n627) );
  XNOR2_X1 U916 ( .A(n143), .B(\fence_regs_cta_id_in[13><3] ), .ZN(n626) );
  NAND2_X1 U917 ( .A1(n528), .A2(warps_per_block_in[2]), .ZN(n625) );
  INV_X1 U918 ( .A(n480), .ZN(n528) );
  NAND2_X1 U919 ( .A1(warps_per_block_in[3]), .A2(warps_per_block_in[1]), .ZN(
        n480) );
  AOI21_X1 U920 ( .B1(n615), .B2(n630), .A(n472), .ZN(cta_id_mask_rev[12]) );
  NAND4_X1 U921 ( .A1(n631), .A2(n632), .A3(n633), .A4(n634), .ZN(n472) );
  XNOR2_X1 U922 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[12><0] ), .ZN(
        n634) );
  XNOR2_X1 U923 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[12><1] ), .ZN(
        n633) );
  XNOR2_X1 U924 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[12><2] ), .ZN(
        n632) );
  XNOR2_X1 U925 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[12><3] ), .ZN(
        n631) );
  NAND2_X1 U926 ( .A1(n546), .A2(warps_per_block_in[2]), .ZN(n630) );
  INV_X1 U927 ( .A(n485), .ZN(n546) );
  NAND2_X1 U928 ( .A1(warps_per_block_in[3]), .A2(n512), .ZN(n485) );
  INV_X1 U929 ( .A(n635), .ZN(n512) );
  NOR2_X1 U930 ( .A1(n479), .A2(n474), .ZN(cta_id_mask_rev[11]) );
  NAND4_X1 U931 ( .A1(n636), .A2(n637), .A3(n638), .A4(n639), .ZN(n474) );
  XNOR2_X1 U932 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[11><0] ), .ZN(
        n639) );
  XNOR2_X1 U933 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[11><1] ), .ZN(
        n638) );
  XNOR2_X1 U934 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[11><2] ), .ZN(
        n637) );
  XNOR2_X1 U935 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[11><3] ), .ZN(
        n636) );
  AOI21_X1 U936 ( .B1(warps_per_block_in[3]), .B2(warps_per_block_in[2]), .A(
        n640), .ZN(n479) );
  AOI21_X1 U937 ( .B1(n615), .B2(n641), .A(n476), .ZN(cta_id_mask_rev[10]) );
  NAND4_X1 U938 ( .A1(n642), .A2(n643), .A3(n644), .A4(n645), .ZN(n476) );
  XNOR2_X1 U939 ( .A(cta_id_in[0]), .B(\fence_regs_cta_id_in[10><0] ), .ZN(
        n645) );
  XNOR2_X1 U940 ( .A(cta_id_in[1]), .B(\fence_regs_cta_id_in[10><1] ), .ZN(
        n644) );
  XNOR2_X1 U941 ( .A(cta_id_in[2]), .B(\fence_regs_cta_id_in[10><2] ), .ZN(
        n643) );
  XNOR2_X1 U942 ( .A(cta_id_in[3]), .B(\fence_regs_cta_id_in[10><3] ), .ZN(
        n642) );
  NAND2_X1 U943 ( .A1(warps_per_block_in[3]), .A2(n557), .ZN(n641) );
  INV_X1 U944 ( .A(n530), .ZN(n557) );
  NOR2_X1 U945 ( .A1(warps_per_block_in[2]), .A2(n500), .ZN(n530) );
  AND2_X1 U946 ( .A1(warps_per_block_in[0]), .A2(warps_per_block_in[1]), .ZN(
        n500) );
  AOI21_X1 U947 ( .B1(n635), .B2(n513), .A(n478), .ZN(cta_id_mask_rev[0]) );
  NAND4_X1 U948 ( .A1(n646), .A2(n647), .A3(n648), .A4(n649), .ZN(n478) );
  XNOR2_X1 U949 ( .A(n137), .B(\fence_regs_cta_id_in[0><0] ), .ZN(n649) );
  XNOR2_X1 U950 ( .A(n139), .B(\fence_regs_cta_id_in[0><1] ), .ZN(n648) );
  XNOR2_X1 U951 ( .A(n141), .B(\fence_regs_cta_id_in[0><2] ), .ZN(n647) );
  XNOR2_X1 U952 ( .A(n143), .B(\fence_regs_cta_id_in[0><3] ), .ZN(n646) );
  NOR2_X1 U953 ( .A1(n501), .A2(warps_per_block_in[2]), .ZN(n513) );
  INV_X1 U954 ( .A(n490), .ZN(n501) );
  NOR2_X1 U955 ( .A1(n640), .A2(warps_per_block_in[3]), .ZN(n490) );
  INV_X1 U956 ( .A(n615), .ZN(n640) );
  NOR2_X1 U957 ( .A1(n540), .A2(warps_per_block_in[4]), .ZN(n615) );
  NAND4_X1 U958 ( .A1(n142), .A2(n144), .A3(n140), .A4(n650), .ZN(n540) );
  NOR2_X1 U959 ( .A1(cta_id_in[0]), .A2(N1190), .ZN(n650) );
  NOR2_X1 U960 ( .A1(warps_per_block_in[1]), .A2(warps_per_block_in[0]), .ZN(
        n635) );
endmodule
