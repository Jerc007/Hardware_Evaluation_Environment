/* -------------------------------------------------------------------------
-- Company:          
-- Engineer:         
-- 
-- Create Date:      
-- Module Name:      warp_scheduler - post_syn. 
-- Project Name:     GPGPU
-- Target Devices: 
-- Tool versions:    
-- Description: 
--
----------------------------------------------------------------------------
---------------------------------------------------------------------------- */

module warp_scheduler_SHMEM_ADDR_SIZE14_DW01_cmp6_1 ( A, B, TC, LT, GT, EQ, LE, 
        GE, NE );
  input [31:0] A;
  input [31:0] B;
  input TC;
  output LT, GT, EQ, LE, GE, NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;

  INV_X1 U1 ( .A(A[1]), .ZN(n2) );
  INV_X1 U2 ( .A(A[0]), .ZN(n3) );
  INV_X1 U3 ( .A(B[1]), .ZN(n1) );
  NOR4_X1 U4 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(EQ) );
  NAND4_X1 U5 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .ZN(n7) );
  XNOR2_X1 U6 ( .A(B[3]), .B(A[3]), .ZN(n11) );
  XNOR2_X1 U7 ( .A(B[4]), .B(A[4]), .ZN(n10) );
  XNOR2_X1 U8 ( .A(B[5]), .B(A[5]), .ZN(n9) );
  XNOR2_X1 U9 ( .A(B[6]), .B(A[6]), .ZN(n8) );
  NAND4_X1 U10 ( .A1(n12), .A2(n13), .A3(n14), .A4(n15), .ZN(n6) );
  OAI22_X1 U11 ( .A1(n16), .A2(n2), .B1(B[1]), .B2(n16), .ZN(n15) );
  AND2_X1 U12 ( .A1(B[0]), .A2(n3), .ZN(n16) );
  OAI22_X1 U13 ( .A1(A[1]), .A2(n17), .B1(n17), .B2(n1), .ZN(n14) );
  NOR2_X1 U14 ( .A1(n3), .A2(B[0]), .ZN(n17) );
  XNOR2_X1 U15 ( .A(B[31]), .B(A[31]), .ZN(n13) );
  XNOR2_X1 U16 ( .A(B[2]), .B(A[2]), .ZN(n12) );
  NAND2_X1 U17 ( .A1(n18), .A2(n19), .ZN(n5) );
  NOR4_X1 U18 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .ZN(n19) );
  XOR2_X1 U19 ( .A(B[10]), .B(A[10]), .Z(n23) );
  XOR2_X1 U20 ( .A(B[9]), .B(A[9]), .Z(n22) );
  XOR2_X1 U21 ( .A(B[8]), .B(A[8]), .Z(n21) );
  XOR2_X1 U22 ( .A(B[7]), .B(A[7]), .Z(n20) );
  NOR4_X1 U23 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(n18) );
  XOR2_X1 U24 ( .A(B[14]), .B(A[14]), .Z(n27) );
  XOR2_X1 U25 ( .A(B[13]), .B(A[13]), .Z(n26) );
  XOR2_X1 U26 ( .A(B[12]), .B(A[12]), .Z(n25) );
  XOR2_X1 U27 ( .A(B[11]), .B(A[11]), .Z(n24) );
  NAND4_X1 U28 ( .A1(n28), .A2(n29), .A3(n30), .A4(n31), .ZN(n4) );
  NOR4_X1 U29 ( .A1(n32), .A2(n33), .A3(n34), .A4(n35), .ZN(n31) );
  XOR2_X1 U30 ( .A(B[18]), .B(A[18]), .Z(n35) );
  XOR2_X1 U31 ( .A(B[17]), .B(A[17]), .Z(n34) );
  XOR2_X1 U32 ( .A(B[16]), .B(A[16]), .Z(n33) );
  XOR2_X1 U33 ( .A(B[15]), .B(A[15]), .Z(n32) );
  NOR4_X1 U34 ( .A1(n36), .A2(n37), .A3(n38), .A4(n39), .ZN(n30) );
  XOR2_X1 U35 ( .A(B[22]), .B(A[22]), .Z(n39) );
  XOR2_X1 U36 ( .A(B[21]), .B(A[21]), .Z(n38) );
  XOR2_X1 U37 ( .A(B[20]), .B(A[20]), .Z(n37) );
  XOR2_X1 U38 ( .A(B[19]), .B(A[19]), .Z(n36) );
  NOR4_X1 U39 ( .A1(n40), .A2(n41), .A3(n42), .A4(n43), .ZN(n29) );
  XOR2_X1 U40 ( .A(B[26]), .B(A[26]), .Z(n43) );
  XOR2_X1 U41 ( .A(B[25]), .B(A[25]), .Z(n42) );
  XOR2_X1 U42 ( .A(B[24]), .B(A[24]), .Z(n41) );
  XOR2_X1 U43 ( .A(B[23]), .B(A[23]), .Z(n40) );
  NOR4_X1 U44 ( .A1(n44), .A2(n45), .A3(n46), .A4(n47), .ZN(n28) );
  XOR2_X1 U45 ( .A(B[30]), .B(A[30]), .Z(n47) );
  XOR2_X1 U46 ( .A(B[29]), .B(A[29]), .Z(n46) );
  XOR2_X1 U47 ( .A(B[28]), .B(A[28]), .Z(n45) );
  XOR2_X1 U48 ( .A(B[27]), .B(A[27]), .Z(n44) );
endmodule



module warp_scheduler ( clk_in, host_reset, reset, 
        pipeline_stall_in, num_blocks_in, num_warps_in, gprs_size_in, 
        warps_done_mask_in, warp_pool_addr_out, warp_pool_wr_en_out, 
        warp_pool_wr_data_out, warp_pool_rd_data_in, warp_state_addr_out, 
        warp_state_wr_en_out, warp_state_wr_data_out, warp_state_rd_data_in, 
        program_cntr_out, warp_id_out, warp_lane_id_out, cta_id_out, 
        initial_mask_out, current_mask_out, shmem_base_addr_out, gprs_size_out, 
        gprs_base_addr_out, done, pipeline_warpunit_done, fetch_en );
  input [3:0] num_blocks_in;
  input [4:0] num_warps_in;
  input [8:0] gprs_size_in;
  input [31:0] warps_done_mask_in;
  output [4:0] warp_pool_addr_out;
  output [127:0] warp_pool_wr_data_out;
  input [127:0] warp_pool_rd_data_in;
  output [4:0] warp_state_addr_out;
  output [1:0] warp_state_wr_data_out;
  input [1:0] warp_state_rd_data_in;
  output [31:0] program_cntr_out;
  output [4:0] warp_id_out;
  output [1:0] warp_lane_id_out;
  output [3:0] cta_id_out;
  output [31:0] initial_mask_out;
  output [31:0] current_mask_out;
  output [13:0] shmem_base_addr_out;
  output [8:0] gprs_size_out;
  output [8:0] gprs_base_addr_out;
  input clk_in, host_reset, reset, pipeline_stall_in;
  output warp_pool_wr_en_out, warp_state_wr_en_out, done,
         pipeline_warpunit_done, fetch_en;
  wire   N52, N63, N64, N66, N67, N70, N71, N72, N73, N94, N321, N322, N323,
         N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334,
         N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345,
         N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356,
         N357, N358, N359, N360, N362, N364, N365, N366, N367, N368, N369,
         N370, N371, N372, N373, N375, N376, N377, N378, N379, N380, N381,
         N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392,
         N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403,
         N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414,
         N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425,
         N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436,
         N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447,
         N448, N449, N450, N451, N452, N453, N454, N455, n161, n166, n167,
         n168, n169, n170, n177, n178, n179, n180, n181, n182, n183, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         \r149/carry[4] , \r149/carry[3] , \r149/carry[2] , n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n162, n163, n164, n165, n171,
         n172, n173, n174, n175, n176, n184, n185, n186, n187, n212, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649;
  wire   [1:0] warp_lane_cnt;
  wire   [4:0] warp_id_cnt;
  wire   [2:0] warp_scheduler_next_state;
  wire   [2:0] warp_scheduler_state_machine;
  wire   [31:0] warps_done_mask;
  assign warp_pool_wr_en_out = 1'b0;
  assign warp_state_wr_data_out[1] = 1'b0;
  assign N321 = warp_pool_rd_data_in[110];
  assign N322 = warp_pool_rd_data_in[111];
  assign N323 = warp_pool_rd_data_in[112];
  assign N324 = warp_pool_rd_data_in[113];
  assign N325 = warp_pool_rd_data_in[114];
  assign N326 = warp_pool_rd_data_in[115];
  assign N327 = warp_pool_rd_data_in[116];
  assign N328 = warp_pool_rd_data_in[117];
  assign N329 = warp_pool_rd_data_in[118];
  assign N330 = warp_pool_rd_data_in[119];
  assign N331 = warp_pool_rd_data_in[120];
  assign N332 = warp_pool_rd_data_in[121];
  assign N333 = warp_pool_rd_data_in[122];
  assign N334 = warp_pool_rd_data_in[123];
  assign N335 = warp_pool_rd_data_in[106];
  assign N336 = warp_pool_rd_data_in[107];
  assign N337 = warp_pool_rd_data_in[108];
  assign N338 = warp_pool_rd_data_in[109];
  assign N339 = warp_pool_rd_data_in[97];
  assign N340 = warp_pool_rd_data_in[98];
  assign N341 = warp_pool_rd_data_in[99];
  assign N342 = warp_pool_rd_data_in[100];
  assign N343 = warp_pool_rd_data_in[101];
  assign N344 = warp_pool_rd_data_in[102];
  assign N345 = warp_pool_rd_data_in[103];
  assign N346 = warp_pool_rd_data_in[104];
  assign N347 = warp_pool_rd_data_in[105];
  assign N348 = warp_pool_rd_data_in[32];
  assign N349 = warp_pool_rd_data_in[33];
  assign N350 = warp_pool_rd_data_in[34];
  assign N351 = warp_pool_rd_data_in[35];
  assign N352 = warp_pool_rd_data_in[36];
  assign N353 = warp_pool_rd_data_in[37];
  assign N354 = warp_pool_rd_data_in[38];
  assign N355 = warp_pool_rd_data_in[39];
  assign N356 = warp_pool_rd_data_in[40];
  assign N357 = warp_pool_rd_data_in[41];
  assign N358 = warp_pool_rd_data_in[42];
  assign N359 = warp_pool_rd_data_in[43];
  assign N360 = warp_pool_rd_data_in[44];
  assign N362 = warp_pool_rd_data_in[45];
  assign N364 = warp_pool_rd_data_in[46];
  assign N365 = warp_pool_rd_data_in[47];
  assign N366 = warp_pool_rd_data_in[48];
  assign N367 = warp_pool_rd_data_in[49];
  assign N368 = warp_pool_rd_data_in[50];
  assign N369 = warp_pool_rd_data_in[51];
  assign N370 = warp_pool_rd_data_in[52];
  assign N371 = warp_pool_rd_data_in[53];
  assign N372 = warp_pool_rd_data_in[54];
  assign N373 = warp_pool_rd_data_in[55];
  assign N375 = warp_pool_rd_data_in[56];
  assign N376 = warp_pool_rd_data_in[57];
  assign N377 = warp_pool_rd_data_in[58];
  assign N378 = warp_pool_rd_data_in[59];
  assign N379 = warp_pool_rd_data_in[60];
  assign N380 = warp_pool_rd_data_in[61];
  assign N381 = warp_pool_rd_data_in[62];
  assign N382 = warp_pool_rd_data_in[63];
  assign N383 = warp_pool_rd_data_in[0];
  assign N384 = warp_pool_rd_data_in[1];
  assign N385 = warp_pool_rd_data_in[2];
  assign N386 = warp_pool_rd_data_in[3];
  assign N387 = warp_pool_rd_data_in[4];
  assign N388 = warp_pool_rd_data_in[5];
  assign N389 = warp_pool_rd_data_in[6];
  assign N390 = warp_pool_rd_data_in[7];
  assign N391 = warp_pool_rd_data_in[8];
  assign N392 = warp_pool_rd_data_in[9];
  assign N393 = warp_pool_rd_data_in[10];
  assign N394 = warp_pool_rd_data_in[11];
  assign N395 = warp_pool_rd_data_in[12];
  assign N396 = warp_pool_rd_data_in[13];
  assign N397 = warp_pool_rd_data_in[14];
  assign N398 = warp_pool_rd_data_in[15];
  assign N399 = warp_pool_rd_data_in[16];
  assign N400 = warp_pool_rd_data_in[17];
  assign N401 = warp_pool_rd_data_in[18];
  assign N402 = warp_pool_rd_data_in[19];
  assign N403 = warp_pool_rd_data_in[20];
  assign N404 = warp_pool_rd_data_in[21];
  assign N405 = warp_pool_rd_data_in[22];
  assign N406 = warp_pool_rd_data_in[23];
  assign N407 = warp_pool_rd_data_in[24];
  assign N408 = warp_pool_rd_data_in[25];
  assign N409 = warp_pool_rd_data_in[26];
  assign N410 = warp_pool_rd_data_in[27];
  assign N411 = warp_pool_rd_data_in[28];
  assign N412 = warp_pool_rd_data_in[29];
  assign N413 = warp_pool_rd_data_in[30];
  assign N414 = warp_pool_rd_data_in[31];
  assign N415 = warp_pool_rd_data_in[64];
  assign N416 = warp_pool_rd_data_in[65];
  assign N417 = warp_pool_rd_data_in[66];
  assign N418 = warp_pool_rd_data_in[67];
  assign N419 = warp_pool_rd_data_in[68];
  assign N420 = warp_pool_rd_data_in[69];
  assign N421 = warp_pool_rd_data_in[70];
  assign N422 = warp_pool_rd_data_in[71];
  assign N423 = warp_pool_rd_data_in[72];
  assign N424 = warp_pool_rd_data_in[73];
  assign N425 = warp_pool_rd_data_in[74];
  assign N426 = warp_pool_rd_data_in[75];
  assign N427 = warp_pool_rd_data_in[76];
  assign N428 = warp_pool_rd_data_in[77];
  assign N429 = warp_pool_rd_data_in[78];
  assign N430 = warp_pool_rd_data_in[79];
  assign N431 = warp_pool_rd_data_in[80];
  assign N432 = warp_pool_rd_data_in[81];
  assign N433 = warp_pool_rd_data_in[82];
  assign N434 = warp_pool_rd_data_in[83];
  assign N435 = warp_pool_rd_data_in[84];
  assign N436 = warp_pool_rd_data_in[85];
  assign N437 = warp_pool_rd_data_in[86];
  assign N438 = warp_pool_rd_data_in[87];
  assign N439 = warp_pool_rd_data_in[88];
  assign N440 = warp_pool_rd_data_in[89];
  assign N441 = warp_pool_rd_data_in[90];
  assign N442 = warp_pool_rd_data_in[91];
  assign N443 = warp_pool_rd_data_in[92];
  assign N444 = warp_pool_rd_data_in[93];
  assign N445 = warp_pool_rd_data_in[94];
  assign N446 = warp_pool_rd_data_in[95];
  assign N447 = gprs_size_in[0];
  assign N448 = gprs_size_in[1];
  assign N449 = gprs_size_in[2];
  assign N450 = gprs_size_in[3];
  assign N451 = gprs_size_in[4];
  assign N452 = gprs_size_in[5];
  assign N453 = gprs_size_in[6];
  assign N454 = gprs_size_in[7];
  assign N455 = gprs_size_in[8];
  assign warp_pool_wr_data_out[127] = 1'b0;
  assign warp_pool_wr_data_out[126] = 1'b0;
  assign warp_pool_wr_data_out[125] = 1'b0;
  assign warp_pool_wr_data_out[124] = 1'b0;
  assign warp_pool_wr_data_out[123] = 1'b0;
  assign warp_pool_wr_data_out[122] = 1'b0;
  assign warp_pool_wr_data_out[121] = 1'b0;
  assign warp_pool_wr_data_out[120] = 1'b0;
  assign warp_pool_wr_data_out[119] = 1'b0;
  assign warp_pool_wr_data_out[118] = 1'b0;
  assign warp_pool_wr_data_out[117] = 1'b0;
  assign warp_pool_wr_data_out[116] = 1'b0;
  assign warp_pool_wr_data_out[115] = 1'b0;
  assign warp_pool_wr_data_out[114] = 1'b0;
  assign warp_pool_wr_data_out[113] = 1'b0;
  assign warp_pool_wr_data_out[112] = 1'b0;
  assign warp_pool_wr_data_out[111] = 1'b0;
  assign warp_pool_wr_data_out[110] = 1'b0;
  assign warp_pool_wr_data_out[109] = 1'b0;
  assign warp_pool_wr_data_out[108] = 1'b0;
  assign warp_pool_wr_data_out[107] = 1'b0;
  assign warp_pool_wr_data_out[106] = 1'b0;
  assign warp_pool_wr_data_out[105] = 1'b0;
  assign warp_pool_wr_data_out[104] = 1'b0;
  assign warp_pool_wr_data_out[103] = 1'b0;
  assign warp_pool_wr_data_out[102] = 1'b0;
  assign warp_pool_wr_data_out[101] = 1'b0;
  assign warp_pool_wr_data_out[100] = 1'b0;
  assign warp_pool_wr_data_out[99] = 1'b0;
  assign warp_pool_wr_data_out[98] = 1'b0;
  assign warp_pool_wr_data_out[97] = 1'b0;
  assign warp_pool_wr_data_out[96] = 1'b0;
  assign warp_pool_wr_data_out[95] = 1'b0;
  assign warp_pool_wr_data_out[94] = 1'b0;
  assign warp_pool_wr_data_out[93] = 1'b0;
  assign warp_pool_wr_data_out[92] = 1'b0;
  assign warp_pool_wr_data_out[91] = 1'b0;
  assign warp_pool_wr_data_out[90] = 1'b0;
  assign warp_pool_wr_data_out[89] = 1'b0;
  assign warp_pool_wr_data_out[88] = 1'b0;
  assign warp_pool_wr_data_out[87] = 1'b0;
  assign warp_pool_wr_data_out[86] = 1'b0;
  assign warp_pool_wr_data_out[85] = 1'b0;
  assign warp_pool_wr_data_out[84] = 1'b0;
  assign warp_pool_wr_data_out[83] = 1'b0;
  assign warp_pool_wr_data_out[82] = 1'b0;
  assign warp_pool_wr_data_out[81] = 1'b0;
  assign warp_pool_wr_data_out[80] = 1'b0;
  assign warp_pool_wr_data_out[79] = 1'b0;
  assign warp_pool_wr_data_out[78] = 1'b0;
  assign warp_pool_wr_data_out[77] = 1'b0;
  assign warp_pool_wr_data_out[76] = 1'b0;
  assign warp_pool_wr_data_out[75] = 1'b0;
  assign warp_pool_wr_data_out[74] = 1'b0;
  assign warp_pool_wr_data_out[73] = 1'b0;
  assign warp_pool_wr_data_out[72] = 1'b0;
  assign warp_pool_wr_data_out[71] = 1'b0;
  assign warp_pool_wr_data_out[70] = 1'b0;
  assign warp_pool_wr_data_out[69] = 1'b0;
  assign warp_pool_wr_data_out[68] = 1'b0;
  assign warp_pool_wr_data_out[67] = 1'b0;
  assign warp_pool_wr_data_out[66] = 1'b0;
  assign warp_pool_wr_data_out[65] = 1'b0;
  assign warp_pool_wr_data_out[64] = 1'b0;
  assign warp_pool_wr_data_out[63] = 1'b0;
  assign warp_pool_wr_data_out[62] = 1'b0;
  assign warp_pool_wr_data_out[61] = 1'b0;
  assign warp_pool_wr_data_out[60] = 1'b0;
  assign warp_pool_wr_data_out[59] = 1'b0;
  assign warp_pool_wr_data_out[58] = 1'b0;
  assign warp_pool_wr_data_out[57] = 1'b0;
  assign warp_pool_wr_data_out[56] = 1'b0;
  assign warp_pool_wr_data_out[55] = 1'b0;
  assign warp_pool_wr_data_out[54] = 1'b0;
  assign warp_pool_wr_data_out[53] = 1'b0;
  assign warp_pool_wr_data_out[52] = 1'b0;
  assign warp_pool_wr_data_out[51] = 1'b0;
  assign warp_pool_wr_data_out[50] = 1'b0;
  assign warp_pool_wr_data_out[49] = 1'b0;
  assign warp_pool_wr_data_out[48] = 1'b0;
  assign warp_pool_wr_data_out[47] = 1'b0;
  assign warp_pool_wr_data_out[46] = 1'b0;
  assign warp_pool_wr_data_out[45] = 1'b0;
  assign warp_pool_wr_data_out[44] = 1'b0;
  assign warp_pool_wr_data_out[43] = 1'b0;
  assign warp_pool_wr_data_out[42] = 1'b0;
  assign warp_pool_wr_data_out[41] = 1'b0;
  assign warp_pool_wr_data_out[40] = 1'b0;
  assign warp_pool_wr_data_out[39] = 1'b0;
  assign warp_pool_wr_data_out[38] = 1'b0;
  assign warp_pool_wr_data_out[37] = 1'b0;
  assign warp_pool_wr_data_out[36] = 1'b0;
  assign warp_pool_wr_data_out[35] = 1'b0;
  assign warp_pool_wr_data_out[34] = 1'b0;
  assign warp_pool_wr_data_out[33] = 1'b0;
  assign warp_pool_wr_data_out[32] = 1'b0;
  assign warp_pool_wr_data_out[31] = 1'b0;
  assign warp_pool_wr_data_out[30] = 1'b0;
  assign warp_pool_wr_data_out[29] = 1'b0;
  assign warp_pool_wr_data_out[28] = 1'b0;
  assign warp_pool_wr_data_out[27] = 1'b0;
  assign warp_pool_wr_data_out[26] = 1'b0;
  assign warp_pool_wr_data_out[25] = 1'b0;
  assign warp_pool_wr_data_out[24] = 1'b0;
  assign warp_pool_wr_data_out[23] = 1'b0;
  assign warp_pool_wr_data_out[22] = 1'b0;
  assign warp_pool_wr_data_out[21] = 1'b0;
  assign warp_pool_wr_data_out[20] = 1'b0;
  assign warp_pool_wr_data_out[19] = 1'b0;
  assign warp_pool_wr_data_out[18] = 1'b0;
  assign warp_pool_wr_data_out[17] = 1'b0;
  assign warp_pool_wr_data_out[16] = 1'b0;
  assign warp_pool_wr_data_out[15] = 1'b0;
  assign warp_pool_wr_data_out[14] = 1'b0;
  assign warp_pool_wr_data_out[13] = 1'b0;
  assign warp_pool_wr_data_out[12] = 1'b0;
  assign warp_pool_wr_data_out[11] = 1'b0;
  assign warp_pool_wr_data_out[10] = 1'b0;
  assign warp_pool_wr_data_out[9] = 1'b0;
  assign warp_pool_wr_data_out[8] = 1'b0;
  assign warp_pool_wr_data_out[7] = 1'b0;
  assign warp_pool_wr_data_out[6] = 1'b0;
  assign warp_pool_wr_data_out[5] = 1'b0;
  assign warp_pool_wr_data_out[4] = 1'b0;
  assign warp_pool_wr_data_out[3] = 1'b0;
  assign warp_pool_wr_data_out[2] = 1'b0;
  assign warp_pool_wr_data_out[1] = 1'b0;
  assign warp_pool_wr_data_out[0] = 1'b0;

  DFFR_X1 \warp_scheduler_next_state_reg[0]  ( .D(n430), .CK(clk_in), .RN(n150), .Q(warp_scheduler_next_state[0]), .QN(n183) );
  DFFR_X1 \warp_scheduler_state_machine_reg[0]  ( .D(n428), .CK(clk_in), .RN(
        n150), .Q(warp_scheduler_state_machine[0]), .QN(n167) );
  DFFR_X1 \warp_lane_cnt_reg[1]  ( .D(n425), .CK(clk_in), .RN(n150), .Q(
        warp_lane_cnt[1]), .QN(n168) );
  DFFR_X1 \warp_scheduler_next_state_reg[2]  ( .D(n421), .CK(clk_in), .RN(n150), .Q(warp_scheduler_next_state[2]), .QN(n181) );
  DFFR_X1 \warp_scheduler_state_machine_reg[2]  ( .D(n429), .CK(clk_in), .RN(
        n150), .Q(warp_scheduler_state_machine[2]), .QN(n161) );
  DFFR_X1 \initial_mask_out_reg[12]  ( .D(n500), .CK(clk_in), .RN(n150), .Q(
        initial_mask_out[12]) );
  DFFR_X1 \initial_mask_out_reg[11]  ( .D(n501), .CK(clk_in), .RN(n150), .Q(
        initial_mask_out[11]) );
  DFFR_X1 \initial_mask_out_reg[10]  ( .D(n502), .CK(clk_in), .RN(n150), .Q(
        initial_mask_out[10]) );
  DFFR_X1 \initial_mask_out_reg[9]  ( .D(n503), .CK(clk_in), .RN(n150), .Q(
        initial_mask_out[9]) );
  DFFR_X1 \initial_mask_out_reg[8]  ( .D(n504), .CK(clk_in), .RN(n150), .Q(
        initial_mask_out[8]) );
  DFFR_X1 \initial_mask_out_reg[7]  ( .D(n505), .CK(clk_in), .RN(n150), .Q(
        initial_mask_out[7]) );
  DFFR_X1 \initial_mask_out_reg[6]  ( .D(n506), .CK(clk_in), .RN(n149), .Q(
        initial_mask_out[6]) );
  DFFR_X1 \initial_mask_out_reg[5]  ( .D(n507), .CK(clk_in), .RN(n149), .Q(
        initial_mask_out[5]) );
  DFFR_X1 \initial_mask_out_reg[4]  ( .D(n508), .CK(clk_in), .RN(n149), .Q(
        initial_mask_out[4]) );
  DFFR_X1 \initial_mask_out_reg[3]  ( .D(n509), .CK(clk_in), .RN(n149), .Q(
        initial_mask_out[3]) );
  DFFR_X1 \initial_mask_out_reg[2]  ( .D(n510), .CK(clk_in), .RN(n149), .Q(
        initial_mask_out[2]) );
  DFFR_X1 \initial_mask_out_reg[1]  ( .D(n511), .CK(clk_in), .RN(n149), .Q(
        initial_mask_out[1]) );
  DFFR_X1 \initial_mask_out_reg[0]  ( .D(n512), .CK(clk_in), .RN(n149), .Q(
        initial_mask_out[0]) );
  DFFR_X1 \gprs_base_addr_out_reg[8]  ( .D(n513), .CK(clk_in), .RN(n149), .Q(
        gprs_base_addr_out[8]) );
  DFFR_X1 \gprs_base_addr_out_reg[7]  ( .D(n514), .CK(clk_in), .RN(n149), .Q(
        gprs_base_addr_out[7]) );
  DFFR_X1 \gprs_base_addr_out_reg[6]  ( .D(n515), .CK(clk_in), .RN(n149), .Q(
        gprs_base_addr_out[6]) );
  DFFR_X1 \gprs_base_addr_out_reg[5]  ( .D(n516), .CK(clk_in), .RN(n149), .Q(
        gprs_base_addr_out[5]) );
  DFFR_X1 \gprs_base_addr_out_reg[4]  ( .D(n517), .CK(clk_in), .RN(n149), .Q(
        gprs_base_addr_out[4]) );
  DFFR_X1 \gprs_base_addr_out_reg[3]  ( .D(n518), .CK(clk_in), .RN(n148), .Q(
        gprs_base_addr_out[3]) );
  DFFR_X1 \gprs_base_addr_out_reg[2]  ( .D(n519), .CK(clk_in), .RN(n148), .Q(
        gprs_base_addr_out[2]) );
  DFFR_X1 \gprs_base_addr_out_reg[1]  ( .D(n520), .CK(clk_in), .RN(n148), .Q(
        gprs_base_addr_out[1]) );
  DFFR_X1 \gprs_base_addr_out_reg[0]  ( .D(n521), .CK(clk_in), .RN(n148), .Q(
        gprs_base_addr_out[0]) );
  DFFR_X1 \cta_id_out_reg[3]  ( .D(n522), .CK(clk_in), .RN(n148), .Q(
        cta_id_out[3]) );
  DFFR_X1 \cta_id_out_reg[2]  ( .D(n523), .CK(clk_in), .RN(n148), .Q(
        cta_id_out[2]) );
  DFFR_X1 \cta_id_out_reg[1]  ( .D(n524), .CK(clk_in), .RN(n148), .Q(
        cta_id_out[1]) );
  DFFR_X1 \cta_id_out_reg[0]  ( .D(n525), .CK(clk_in), .RN(n148), .Q(
        cta_id_out[0]) );
  DFFR_X1 \shmem_base_addr_out_reg[13]  ( .D(n526), .CK(clk_in), .RN(n148), 
        .Q(shmem_base_addr_out[13]) );
  DFFR_X1 \shmem_base_addr_out_reg[12]  ( .D(n527), .CK(clk_in), .RN(n148), 
        .Q(shmem_base_addr_out[12]) );
  DFFR_X1 \shmem_base_addr_out_reg[11]  ( .D(n528), .CK(clk_in), .RN(n148), 
        .Q(shmem_base_addr_out[11]) );
  DFFR_X1 \shmem_base_addr_out_reg[10]  ( .D(n529), .CK(clk_in), .RN(n148), 
        .Q(shmem_base_addr_out[10]) );
  DFFR_X1 \shmem_base_addr_out_reg[9]  ( .D(n530), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[9]) );
  DFFR_X1 \shmem_base_addr_out_reg[8]  ( .D(n531), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[8]) );
  DFFR_X1 \shmem_base_addr_out_reg[7]  ( .D(n532), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[7]) );
  DFFR_X1 \shmem_base_addr_out_reg[6]  ( .D(n533), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[6]) );
  DFFR_X1 \shmem_base_addr_out_reg[5]  ( .D(n534), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[5]) );
  DFFR_X1 \shmem_base_addr_out_reg[4]  ( .D(n535), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[4]) );
  DFFR_X1 \shmem_base_addr_out_reg[3]  ( .D(n536), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[3]) );
  DFFR_X1 \shmem_base_addr_out_reg[2]  ( .D(n537), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[2]) );
  DFFR_X1 \shmem_base_addr_out_reg[1]  ( .D(n538), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[1]) );
  DFFR_X1 \shmem_base_addr_out_reg[0]  ( .D(n539), .CK(clk_in), .RN(n147), .Q(
        shmem_base_addr_out[0]) );
  DFFR_X1 \gprs_size_out_reg[8]  ( .D(n540), .CK(clk_in), .RN(n147), .Q(
        gprs_size_out[8]) );
  DFFR_X1 \gprs_size_out_reg[7]  ( .D(n541), .CK(clk_in), .RN(n147), .Q(
        gprs_size_out[7]) );
  DFFR_X1 \gprs_size_out_reg[6]  ( .D(n542), .CK(clk_in), .RN(n146), .Q(
        gprs_size_out[6]) );
  DFFR_X1 \gprs_size_out_reg[5]  ( .D(n543), .CK(clk_in), .RN(n146), .Q(
        gprs_size_out[5]) );
  DFFR_X1 \gprs_size_out_reg[4]  ( .D(n544), .CK(clk_in), .RN(n146), .Q(
        gprs_size_out[4]) );
  DFFR_X1 \gprs_size_out_reg[3]  ( .D(n545), .CK(clk_in), .RN(n146), .Q(
        gprs_size_out[3]) );
  DFFR_X1 \gprs_size_out_reg[2]  ( .D(n546), .CK(clk_in), .RN(n146), .Q(
        gprs_size_out[2]) );
  DFFR_X1 \gprs_size_out_reg[1]  ( .D(n547), .CK(clk_in), .RN(n146), .Q(
        gprs_size_out[1]) );
  DFFR_X1 \gprs_size_out_reg[0]  ( .D(n548), .CK(clk_in), .RN(n146), .Q(
        gprs_size_out[0]) );
  DFFR_X1 \program_cntr_out_reg[31]  ( .D(n549), .CK(clk_in), .RN(n146), .Q(
        program_cntr_out[31]) );
  DFFR_X1 \program_cntr_out_reg[30]  ( .D(n550), .CK(clk_in), .RN(n146), .Q(
        program_cntr_out[30]) );
  DFFR_X1 \program_cntr_out_reg[29]  ( .D(n551), .CK(clk_in), .RN(n146), .Q(
        program_cntr_out[29]) );
  DFFR_X1 \program_cntr_out_reg[28]  ( .D(n552), .CK(clk_in), .RN(n146), .Q(
        program_cntr_out[28]) );
  DFFR_X1 \program_cntr_out_reg[27]  ( .D(n553), .CK(clk_in), .RN(n146), .Q(
        program_cntr_out[27]) );
  DFFR_X1 \program_cntr_out_reg[26]  ( .D(n554), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[26]) );
  DFFR_X1 \program_cntr_out_reg[25]  ( .D(n555), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[25]) );
  DFFR_X1 \program_cntr_out_reg[24]  ( .D(n556), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[24]) );
  DFFR_X1 \program_cntr_out_reg[23]  ( .D(n557), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[23]) );
  DFFR_X1 \program_cntr_out_reg[22]  ( .D(n558), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[22]) );
  DFFR_X1 \program_cntr_out_reg[21]  ( .D(n559), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[21]) );
  DFFR_X1 \program_cntr_out_reg[20]  ( .D(n560), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[20]) );
  DFFR_X1 \program_cntr_out_reg[19]  ( .D(n561), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[19]) );
  DFFR_X1 \program_cntr_out_reg[18]  ( .D(n562), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[18]) );
  DFFR_X1 \program_cntr_out_reg[17]  ( .D(n563), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[17]) );
  DFFR_X1 \program_cntr_out_reg[16]  ( .D(n564), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[16]) );
  DFFR_X1 \program_cntr_out_reg[15]  ( .D(n565), .CK(clk_in), .RN(n145), .Q(
        program_cntr_out[15]) );
  DFFR_X1 \program_cntr_out_reg[14]  ( .D(n566), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[14]) );
  DFFR_X1 \program_cntr_out_reg[13]  ( .D(n567), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[13]) );
  DFFR_X1 \program_cntr_out_reg[12]  ( .D(n568), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[12]) );
  DFFR_X1 \program_cntr_out_reg[11]  ( .D(n569), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[11]) );
  DFFR_X1 \program_cntr_out_reg[10]  ( .D(n570), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[10]) );
  DFFR_X1 \program_cntr_out_reg[9]  ( .D(n571), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[9]) );
  DFFR_X1 \program_cntr_out_reg[8]  ( .D(n572), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[8]) );
  DFFR_X1 \program_cntr_out_reg[7]  ( .D(n573), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[7]) );
  DFFR_X1 \program_cntr_out_reg[6]  ( .D(n574), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[6]) );
  DFFR_X1 \program_cntr_out_reg[5]  ( .D(n575), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[5]) );
  DFFR_X1 \program_cntr_out_reg[4]  ( .D(n576), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[4]) );
  DFFR_X1 \program_cntr_out_reg[3]  ( .D(n577), .CK(clk_in), .RN(n144), .Q(
        program_cntr_out[3]) );
  DFFR_X1 \program_cntr_out_reg[2]  ( .D(n578), .CK(clk_in), .RN(n143), .Q(
        program_cntr_out[2]) );
  DFFR_X1 \program_cntr_out_reg[1]  ( .D(n579), .CK(clk_in), .RN(n143), .Q(
        program_cntr_out[1]) );
  DFFR_X1 \program_cntr_out_reg[0]  ( .D(n580), .CK(clk_in), .RN(n143), .Q(
        program_cntr_out[0]) );
  DFFR_X1 \current_mask_out_reg[31]  ( .D(n581), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[31]) );
  DFFR_X1 \current_mask_out_reg[30]  ( .D(n582), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[30]) );
  DFFR_X1 \current_mask_out_reg[29]  ( .D(n583), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[29]) );
  DFFR_X1 \current_mask_out_reg[28]  ( .D(n584), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[28]) );
  DFFR_X1 \current_mask_out_reg[27]  ( .D(n585), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[27]) );
  DFFR_X1 \current_mask_out_reg[26]  ( .D(n586), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[26]) );
  DFFR_X1 \current_mask_out_reg[25]  ( .D(n587), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[25]) );
  DFFR_X1 \current_mask_out_reg[24]  ( .D(n588), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[24]) );
  DFFR_X1 \current_mask_out_reg[23]  ( .D(n589), .CK(clk_in), .RN(n143), .Q(
        current_mask_out[23]) );
  DFFR_X1 \current_mask_out_reg[22]  ( .D(n590), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[22]) );
  DFFR_X1 \current_mask_out_reg[21]  ( .D(n591), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[21]) );
  DFFR_X1 \current_mask_out_reg[20]  ( .D(n592), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[20]) );
  DFFR_X1 \current_mask_out_reg[19]  ( .D(n593), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[19]) );
  DFFR_X1 \current_mask_out_reg[18]  ( .D(n594), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[18]) );
  DFFR_X1 \current_mask_out_reg[17]  ( .D(n595), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[17]) );
  DFFR_X1 \current_mask_out_reg[16]  ( .D(n596), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[16]) );
  DFFR_X1 \current_mask_out_reg[15]  ( .D(n597), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[15]) );
  DFFR_X1 \current_mask_out_reg[14]  ( .D(n598), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[14]) );
  DFFR_X1 \current_mask_out_reg[13]  ( .D(n599), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[13]) );
  DFFR_X1 \current_mask_out_reg[12]  ( .D(n600), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[12]) );
  DFFR_X1 \current_mask_out_reg[11]  ( .D(n601), .CK(clk_in), .RN(n142), .Q(
        current_mask_out[11]) );
  DFFR_X1 \current_mask_out_reg[10]  ( .D(n602), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[10]) );
  DFFR_X1 \current_mask_out_reg[9]  ( .D(n603), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[9]) );
  DFFR_X1 \current_mask_out_reg[8]  ( .D(n604), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[8]) );
  DFFR_X1 \current_mask_out_reg[7]  ( .D(n605), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[7]) );
  DFFR_X1 \current_mask_out_reg[6]  ( .D(n606), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[6]) );
  DFFR_X1 \current_mask_out_reg[5]  ( .D(n607), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[5]) );
  DFFR_X1 \current_mask_out_reg[4]  ( .D(n608), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[4]) );
  DFFR_X1 \current_mask_out_reg[3]  ( .D(n609), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[3]) );
  DFFR_X1 \current_mask_out_reg[2]  ( .D(n610), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[2]) );
  DFFR_X1 \current_mask_out_reg[1]  ( .D(n611), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[1]) );
  DFFR_X1 \current_mask_out_reg[0]  ( .D(n612), .CK(clk_in), .RN(n141), .Q(
        current_mask_out[0]) );
  DFFR_X1 \initial_mask_out_reg[31]  ( .D(n613), .CK(clk_in), .RN(n141), .Q(
        initial_mask_out[31]) );
  DFFR_X1 \initial_mask_out_reg[30]  ( .D(n614), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[30]) );
  DFFR_X1 \initial_mask_out_reg[29]  ( .D(n615), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[29]) );
  DFFR_X1 \initial_mask_out_reg[28]  ( .D(n616), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[28]) );
  DFFR_X1 \initial_mask_out_reg[27]  ( .D(n617), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[27]) );
  DFFR_X1 \initial_mask_out_reg[26]  ( .D(n618), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[26]) );
  DFFR_X1 \initial_mask_out_reg[25]  ( .D(n619), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[25]) );
  DFFR_X1 \initial_mask_out_reg[24]  ( .D(n620), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[24]) );
  DFFR_X1 \initial_mask_out_reg[23]  ( .D(n621), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[23]) );
  DFFR_X1 \initial_mask_out_reg[22]  ( .D(n622), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[22]) );
  DFFR_X1 \initial_mask_out_reg[21]  ( .D(n623), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[21]) );
  DFFR_X1 \initial_mask_out_reg[20]  ( .D(n624), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[20]) );
  DFFR_X1 \initial_mask_out_reg[19]  ( .D(n625), .CK(clk_in), .RN(n140), .Q(
        initial_mask_out[19]) );
  DFFR_X1 \initial_mask_out_reg[18]  ( .D(n626), .CK(clk_in), .RN(n139), .Q(
        initial_mask_out[18]) );
  DFFR_X1 \initial_mask_out_reg[17]  ( .D(n627), .CK(clk_in), .RN(n139), .Q(
        initial_mask_out[17]) );
  DFFR_X1 \initial_mask_out_reg[16]  ( .D(n628), .CK(clk_in), .RN(n139), .Q(
        initial_mask_out[16]) );
  DFFR_X1 \initial_mask_out_reg[15]  ( .D(n629), .CK(clk_in), .RN(n139), .Q(
        initial_mask_out[15]) );
  DFFR_X1 \initial_mask_out_reg[14]  ( .D(n630), .CK(clk_in), .RN(n139), .Q(
        initial_mask_out[14]) );
  DFFR_X1 \initial_mask_out_reg[13]  ( .D(n631), .CK(clk_in), .RN(n139), .Q(
        initial_mask_out[13]) );
  DFFR_X1 \warp_scheduler_next_state_reg[1]  ( .D(n422), .CK(clk_in), .RN(n139), .Q(warp_scheduler_next_state[1]), .QN(n182) );
  DFFR_X1 \warp_scheduler_state_machine_reg[1]  ( .D(n427), .CK(clk_in), .RN(
        n139), .Q(warp_scheduler_state_machine[1]), .QN(n166) );
  DFFR_X1 done_reg ( .D(n638), .CK(clk_in), .RN(n139), .Q(done) );
  DFFR_X1 \warp_state_wr_data_out_reg[0]  ( .D(n419), .CK(clk_in), .RN(n139), 
        .Q(warp_state_wr_data_out[0]) );
  DFFR_X1 warp_state_wr_en_out_reg ( .D(n420), .CK(clk_in), .RN(n139), .Q(
        warp_state_wr_en_out) );
  DFFR_X1 \warp_id_cnt_reg[1]  ( .D(n418), .CK(clk_in), .RN(n139), .Q(
        warp_id_cnt[1]), .QN(n179) );
  DFFR_X1 \warp_id_cnt_reg[4]  ( .D(n414), .CK(clk_in), .RN(n138), .Q(
        warp_id_cnt[4]), .QN(n170) );
  DFFR_X1 \warp_id_cnt_reg[3]  ( .D(n415), .CK(clk_in), .RN(n138), .Q(
        warp_id_cnt[3]), .QN(n177) );
  DFFR_X1 \warp_state_addr_out_reg[3]  ( .D(n405), .CK(clk_in), .RN(n138), .Q(
        warp_state_addr_out[3]) );
  DFFR_X1 \warp_pool_addr_out_reg[3]  ( .D(n410), .CK(clk_in), .RN(n138), .Q(
        warp_pool_addr_out[3]) );
  DFFR_X1 \warp_id_out_reg[3]  ( .D(n494), .CK(clk_in), .RN(n138), .Q(
        warp_id_out[3]) );
  DFFR_X1 \warp_id_cnt_reg[2]  ( .D(n416), .CK(clk_in), .RN(n138), .Q(
        warp_id_cnt[2]), .QN(n178) );
  DFFR_X1 \warp_state_addr_out_reg[2]  ( .D(n406), .CK(clk_in), .RN(n138), .Q(
        warp_state_addr_out[2]) );
  DFFR_X1 \warp_pool_addr_out_reg[2]  ( .D(n411), .CK(clk_in), .RN(n138), .Q(
        warp_pool_addr_out[2]) );
  DFFR_X1 \warp_id_out_reg[2]  ( .D(n495), .CK(clk_in), .RN(n138), .Q(
        warp_id_out[2]) );
  DFFR_X1 \warp_id_cnt_reg[0]  ( .D(n417), .CK(clk_in), .RN(n138), .Q(
        warp_id_cnt[0]), .QN(n180) );
  DFFR_X1 \warp_state_addr_out_reg[0]  ( .D(n408), .CK(clk_in), .RN(n138), .Q(
        warp_state_addr_out[0]) );
  DFFR_X1 \warp_pool_addr_out_reg[0]  ( .D(n413), .CK(clk_in), .RN(n138), .Q(
        warp_pool_addr_out[0]) );
  DFFR_X1 \warp_id_out_reg[0]  ( .D(n496), .CK(clk_in), .RN(n137), .Q(
        warp_id_out[0]) );
  DFFR_X1 \warp_state_addr_out_reg[4]  ( .D(n404), .CK(clk_in), .RN(n137), .Q(
        warp_state_addr_out[4]) );
  DFFR_X1 \warp_pool_addr_out_reg[4]  ( .D(n409), .CK(clk_in), .RN(n137), .Q(
        warp_pool_addr_out[4]) );
  DFFR_X1 \warp_id_out_reg[4]  ( .D(n493), .CK(clk_in), .RN(n137), .Q(
        warp_id_out[4]) );
  DFFR_X1 \warp_state_addr_out_reg[1]  ( .D(n407), .CK(clk_in), .RN(n137), .Q(
        warp_state_addr_out[1]) );
  DFFR_X1 \warp_pool_addr_out_reg[1]  ( .D(n412), .CK(clk_in), .RN(n137), .Q(
        warp_pool_addr_out[1]) );
  DFFR_X1 \warp_id_out_reg[1]  ( .D(n497), .CK(clk_in), .RN(n137), .Q(
        warp_id_out[1]) );
  DFFR_X1 pipeline_warpunit_done_reg ( .D(n426), .CK(clk_in), .RN(n137), .Q(
        pipeline_warpunit_done) );
  DFFR_X1 fetch_en_reg ( .D(n424), .CK(clk_in), .RN(n137), .Q(fetch_en) );
  DFFR_X1 \warp_lane_cnt_reg[0]  ( .D(n423), .CK(clk_in), .RN(n137), .Q(
        warp_lane_cnt[0]), .QN(n169) );
  DFFR_X1 \warp_lane_id_out_reg[0]  ( .D(n498), .CK(clk_in), .RN(n137), .Q(
        warp_lane_id_out[0]) );
  DFFR_X1 \warp_lane_id_out_reg[1]  ( .D(n499), .CK(clk_in), .RN(n137), .Q(
        warp_lane_id_out[1]) );
  NAND2_X1 U382 ( .A1(warp_state_addr_out[4]), .A2(n632), .ZN(n190) );
  NAND2_X1 U383 ( .A1(warp_state_addr_out[3]), .A2(n632), .ZN(n192) );
  NAND2_X1 U384 ( .A1(warp_state_addr_out[2]), .A2(n632), .ZN(n194) );
  NAND2_X1 U385 ( .A1(warp_state_addr_out[1]), .A2(n632), .ZN(n196) );
  NAND2_X1 U386 ( .A1(warp_state_addr_out[0]), .A2(n632), .ZN(n198) );
  NAND2_X1 U387 ( .A1(n202), .A2(n203), .ZN(n199) );
  NAND2_X1 U388 ( .A1(warp_pool_addr_out[4]), .A2(n202), .ZN(n204) );
  NAND2_X1 U389 ( .A1(N73), .A2(n205), .ZN(n189) );
  NAND2_X1 U390 ( .A1(warp_pool_addr_out[3]), .A2(n202), .ZN(n206) );
  NAND2_X1 U391 ( .A1(N72), .A2(n205), .ZN(n191) );
  NAND2_X1 U392 ( .A1(warp_pool_addr_out[2]), .A2(n202), .ZN(n207) );
  NAND2_X1 U393 ( .A1(N71), .A2(n205), .ZN(n193) );
  NAND2_X1 U394 ( .A1(warp_pool_addr_out[1]), .A2(n202), .ZN(n208) );
  NAND2_X1 U395 ( .A1(N70), .A2(n205), .ZN(n195) );
  NAND2_X1 U396 ( .A1(warp_pool_addr_out[0]), .A2(n202), .ZN(n209) );
  NAND2_X1 U397 ( .A1(n180), .A2(n205), .ZN(n197) );
  NAND2_X1 U398 ( .A1(n210), .A2(n221), .ZN(n213) );
  NAND3_X1 U399 ( .A1(n222), .A2(n492), .A3(n223), .ZN(n221) );
  NAND2_X1 U400 ( .A1(n225), .A2(n226), .ZN(n210) );
  NAND2_X1 U401 ( .A1(warp_state_wr_data_out[0]), .A2(n131), .ZN(n228) );
  NAND2_X1 U402 ( .A1(warp_state_wr_en_out), .A2(n229), .ZN(n230) );
  NAND3_X1 U403 ( .A1(n237), .A2(n169), .A3(n239), .ZN(n238) );
  NAND2_X1 U404 ( .A1(fetch_en), .A2(n240), .ZN(n242) );
  NAND3_X1 U405 ( .A1(n239), .A2(n237), .A3(n248), .ZN(n247) );
  NAND2_X1 U406 ( .A1(pipeline_warpunit_done), .A2(n387), .ZN(n388) );
  NAND3_X1 U407 ( .A1(n166), .A2(n161), .A3(n167), .ZN(n392) );
  NAND2_X1 U408 ( .A1(n640), .A2(n231), .ZN(n201) );
  NAND3_X1 U409 ( .A1(warp_scheduler_state_machine[1]), .A2(n167), .A3(
        warp_scheduler_state_machine[2]), .ZN(n231) );
  NAND3_X1 U410 ( .A1(n220), .A2(n232), .A3(n226), .ZN(n235) );
  NAND2_X1 U411 ( .A1(n449), .A2(n403), .ZN(n232) );
  NAND2_X1 U414 ( .A1(n252), .A2(n200), .ZN(n203) );
  warps_done_lut uWarpsDoneLUT ( .clk_in(clk_in), .host_reset(host_reset), 
        .num_warps_in(num_warps_in), .warps_done_mask(warps_done_mask) );
  warp_scheduler_SHMEM_ADDR_SIZE14_DW01_cmp6_1 eq_164 ( .A(warps_done_mask_in), 
        .B(warps_done_mask), .TC(1'b0), .EQ(N52) );
  HA_X1 \r149/U1_1_1  ( .A(warp_id_cnt[1]), .B(warp_id_cnt[0]), .CO(
        \r149/carry[2] ), .S(N70) );
  HA_X1 \r149/U1_1_2  ( .A(warp_id_cnt[2]), .B(\r149/carry[2] ), .CO(
        \r149/carry[3] ), .S(N71) );
  HA_X1 \r149/U1_1_3  ( .A(warp_id_cnt[3]), .B(\r149/carry[3] ), .CO(
        \r149/carry[4] ), .S(N72) );
  NOR3_X1 U133 ( .A1(n167), .A2(warp_scheduler_state_machine[2]), .A3(n166), 
        .ZN(n200) );
  NOR3_X1 U134 ( .A1(warp_scheduler_state_machine[0]), .A2(
        warp_scheduler_state_machine[2]), .A3(n166), .ZN(n244) );
  NOR3_X1 U135 ( .A1(warp_scheduler_state_machine[0]), .A2(
        warp_scheduler_state_machine[1]), .A3(n161), .ZN(n220) );
  AND2_X1 U136 ( .A1(n250), .A2(n203), .ZN(n130) );
  INV_X1 U137 ( .A(n448), .ZN(n154) );
  INV_X1 U138 ( .A(n449), .ZN(n156) );
  INV_X1 U139 ( .A(n447), .ZN(n152) );
  INV_X1 U140 ( .A(n449), .ZN(n157) );
  BUF_X1 U141 ( .A(n450), .Z(n448) );
  BUF_X1 U142 ( .A(n450), .Z(n449) );
  BUF_X1 U143 ( .A(n450), .Z(n447) );
  BUF_X1 U144 ( .A(n451), .Z(n446) );
  BUF_X1 U145 ( .A(n451), .Z(n445) );
  BUF_X1 U146 ( .A(n451), .Z(n444) );
  BUF_X1 U147 ( .A(n452), .Z(n443) );
  BUF_X1 U148 ( .A(n452), .Z(n442) );
  BUF_X1 U149 ( .A(n452), .Z(n441) );
  BUF_X1 U150 ( .A(n453), .Z(n440) );
  BUF_X1 U151 ( .A(n453), .Z(n439) );
  BUF_X1 U152 ( .A(n453), .Z(n438) );
  BUF_X1 U153 ( .A(n454), .Z(n437) );
  BUF_X1 U154 ( .A(n454), .Z(n436) );
  BUF_X1 U155 ( .A(n454), .Z(n435) );
  BUF_X1 U156 ( .A(n455), .Z(n434) );
  BUF_X1 U157 ( .A(n455), .Z(n433) );
  BUF_X1 U158 ( .A(n455), .Z(n432) );
  BUF_X1 U159 ( .A(n456), .Z(n212) );
  BUF_X1 U160 ( .A(n456), .Z(n187) );
  BUF_X1 U161 ( .A(n457), .Z(n186) );
  BUF_X1 U162 ( .A(n457), .Z(n185) );
  BUF_X1 U163 ( .A(n457), .Z(n184) );
  BUF_X1 U164 ( .A(n458), .Z(n176) );
  BUF_X1 U165 ( .A(n458), .Z(n175) );
  BUF_X1 U166 ( .A(n458), .Z(n174) );
  BUF_X1 U167 ( .A(n459), .Z(n173) );
  BUF_X1 U168 ( .A(n459), .Z(n172) );
  BUF_X1 U169 ( .A(n456), .Z(n431) );
  BUF_X1 U170 ( .A(n459), .Z(n171) );
  BUF_X1 U171 ( .A(n460), .Z(n165) );
  BUF_X1 U172 ( .A(n460), .Z(n164) );
  BUF_X1 U173 ( .A(n460), .Z(n163) );
  BUF_X1 U174 ( .A(n461), .Z(n162) );
  BUF_X1 U175 ( .A(n461), .Z(n160) );
  BUF_X1 U176 ( .A(n461), .Z(n159) );
  BUF_X1 U177 ( .A(n462), .Z(n158) );
  BUF_X1 U178 ( .A(n453), .Z(n462) );
  BUF_X1 U179 ( .A(n455), .Z(n457) );
  BUF_X1 U180 ( .A(n453), .Z(n458) );
  BUF_X1 U181 ( .A(n452), .Z(n456) );
  BUF_X1 U182 ( .A(n454), .Z(n459) );
  BUF_X1 U183 ( .A(n453), .Z(n460) );
  BUF_X1 U184 ( .A(n454), .Z(n461) );
  BUF_X1 U185 ( .A(n130), .Z(n450) );
  BUF_X1 U186 ( .A(n130), .Z(n451) );
  BUF_X1 U187 ( .A(n130), .Z(n452) );
  BUF_X1 U188 ( .A(n130), .Z(n453) );
  BUF_X1 U189 ( .A(n130), .Z(n454) );
  BUF_X1 U190 ( .A(n130), .Z(n455) );
  INV_X1 U191 ( .A(n199), .ZN(n632) );
  INV_X1 U192 ( .A(N52), .ZN(n492) );
  NOR2_X1 U193 ( .A1(n492), .A2(n635), .ZN(n397) );
  INV_X1 U194 ( .A(n478), .ZN(n486) );
  AND2_X1 U195 ( .A1(n639), .A2(n210), .ZN(n202) );
  INV_X1 U196 ( .A(n201), .ZN(n639) );
  NOR2_X1 U197 ( .A1(n635), .A2(n648), .ZN(n243) );
  NOR2_X1 U198 ( .A1(n642), .A2(n641), .ZN(n205) );
  AND3_X1 U199 ( .A1(n640), .A2(n203), .A3(n641), .ZN(n131) );
  INV_X1 U200 ( .A(n227), .ZN(n636) );
  INV_X1 U201 ( .A(n223), .ZN(n633) );
  BUF_X1 U202 ( .A(n132), .Z(n134) );
  BUF_X1 U203 ( .A(n132), .Z(n135) );
  BUF_X1 U204 ( .A(n132), .Z(n136) );
  OAI211_X1 U205 ( .C1(n219), .C2(n220), .A(n213), .B(N67), .ZN(n214) );
  INV_X1 U206 ( .A(n220), .ZN(n641) );
  NOR2_X1 U207 ( .A1(n244), .A2(n225), .ZN(n250) );
  INV_X1 U208 ( .A(n398), .ZN(n490) );
  INV_X1 U209 ( .A(n232), .ZN(n491) );
  INV_X1 U210 ( .A(N67), .ZN(n642) );
  INV_X1 U211 ( .A(N66), .ZN(n484) );
  OAI21_X1 U212 ( .B1(n200), .B2(n201), .A(n199), .ZN(n188) );
  OAI21_X1 U213 ( .B1(n249), .B2(n635), .A(n250), .ZN(n237) );
  NOR2_X1 U214 ( .A1(n251), .A2(n252), .ZN(n249) );
  NOR3_X1 U215 ( .A1(n253), .A2(N52), .A3(n254), .ZN(n251) );
  NOR2_X1 U216 ( .A1(n641), .A2(n226), .ZN(n234) );
  NOR2_X1 U217 ( .A1(n244), .A2(n200), .ZN(n227) );
  NOR2_X1 U218 ( .A1(n635), .A2(n254), .ZN(n223) );
  NOR2_X1 U219 ( .A1(n220), .A2(n243), .ZN(n390) );
  NOR2_X1 U220 ( .A1(n647), .A2(n649), .ZN(n253) );
  INV_X1 U221 ( .A(n200), .ZN(n635) );
  INV_X1 U222 ( .A(n244), .ZN(n640) );
  NAND4_X1 U223 ( .A1(n391), .A2(n637), .A3(n640), .A4(n392), .ZN(n245) );
  OR3_X1 U224 ( .A1(n253), .A2(N52), .A3(n635), .ZN(n391) );
  INV_X1 U225 ( .A(n393), .ZN(n637) );
  OR3_X1 U226 ( .A1(n243), .A2(n234), .A3(n244), .ZN(n239) );
  INV_X1 U227 ( .A(n468), .ZN(n485) );
  INV_X1 U228 ( .A(n254), .ZN(n648) );
  NOR2_X1 U229 ( .A1(host_reset), .A2(reset), .ZN(n132) );
  OAI22_X1 U230 ( .A1(warp_state_rd_data_in[1]), .A2(N94), .B1(
        pipeline_stall_in), .B2(n224), .ZN(n222) );
  INV_X1 U231 ( .A(n477), .ZN(n488) );
  NAND4_X1 U232 ( .A1(warp_state_rd_data_in[1]), .A2(n200), .A3(n492), .A4(
        n647), .ZN(n403) );
  OAI211_X1 U233 ( .C1(pipeline_stall_in), .C2(n390), .A(n639), .B(n402), .ZN(
        n398) );
  AOI221_X1 U234 ( .B1(n223), .B2(n649), .C1(warp_scheduler_state_machine[0]), 
        .C2(n166), .A(n397), .ZN(n402) );
  INV_X1 U235 ( .A(n332), .ZN(n577) );
  AOI22_X1 U236 ( .A1(program_cntr_out[3]), .A2(n432), .B1(N418), .B2(n154), 
        .ZN(n332) );
  NOR3_X1 U237 ( .A1(N52), .A2(pipeline_stall_in), .A3(n648), .ZN(n252) );
  NOR2_X1 U238 ( .A1(n641), .A2(pipeline_stall_in), .ZN(n225) );
  XOR2_X1 U239 ( .A(num_warps_in[3]), .B(n465), .Z(n133) );
  OAI221_X1 U240 ( .B1(n491), .B2(n633), .C1(n232), .C2(n182), .A(n235), .ZN(
        n422) );
  OAI22_X1 U241 ( .A1(n180), .A2(n213), .B1(warp_id_cnt[0]), .B2(n214), .ZN(
        n417) );
  OAI22_X1 U242 ( .A1(n178), .A2(n213), .B1(n645), .B2(n214), .ZN(n416) );
  INV_X1 U243 ( .A(N71), .ZN(n645) );
  OAI22_X1 U244 ( .A1(n177), .A2(n213), .B1(n644), .B2(n214), .ZN(n415) );
  INV_X1 U245 ( .A(N72), .ZN(n644) );
  OAI22_X1 U246 ( .A1(n170), .A2(n213), .B1(n643), .B2(n214), .ZN(n414) );
  INV_X1 U247 ( .A(N73), .ZN(n643) );
  OAI22_X1 U248 ( .A1(n179), .A2(n213), .B1(n646), .B2(n214), .ZN(n418) );
  INV_X1 U249 ( .A(N70), .ZN(n646) );
  OAI22_X1 U250 ( .A1(n232), .A2(n181), .B1(n491), .B2(n233), .ZN(n421) );
  NOR2_X1 U251 ( .A1(n234), .A2(n636), .ZN(n233) );
  INV_X1 U252 ( .A(n481), .ZN(n487) );
  AOI21_X1 U253 ( .B1(warp_state_rd_data_in[1]), .B2(n642), .A(n219), .ZN(n224) );
  INV_X1 U254 ( .A(n474), .ZN(n489) );
  OAI21_X1 U255 ( .B1(n232), .B2(n183), .A(n235), .ZN(n430) );
  INV_X1 U256 ( .A(num_warps_in[2]), .ZN(n467) );
  NAND4_X1 U257 ( .A1(n633), .A2(n392), .A3(n231), .A4(n396), .ZN(n427) );
  AOI221_X1 U258 ( .B1(n490), .B2(warp_scheduler_state_machine[1]), .C1(n393), 
        .C2(warp_scheduler_next_state[1]), .A(n397), .ZN(n396) );
  INV_X1 U259 ( .A(n335), .ZN(n580) );
  AOI22_X1 U260 ( .A1(program_cntr_out[0]), .A2(n433), .B1(N415), .B2(n154), 
        .ZN(n335) );
  INV_X1 U261 ( .A(n334), .ZN(n579) );
  AOI22_X1 U262 ( .A1(program_cntr_out[1]), .A2(n432), .B1(N416), .B2(n156), 
        .ZN(n334) );
  INV_X1 U263 ( .A(n333), .ZN(n578) );
  AOI22_X1 U264 ( .A1(program_cntr_out[2]), .A2(n432), .B1(N417), .B2(n151), 
        .ZN(n333) );
  INV_X1 U265 ( .A(n331), .ZN(n576) );
  AOI22_X1 U266 ( .A1(program_cntr_out[4]), .A2(n432), .B1(N419), .B2(n154), 
        .ZN(n331) );
  INV_X1 U267 ( .A(n330), .ZN(n575) );
  AOI22_X1 U268 ( .A1(program_cntr_out[5]), .A2(n431), .B1(N420), .B2(n154), 
        .ZN(n330) );
  INV_X1 U269 ( .A(n329), .ZN(n574) );
  AOI22_X1 U270 ( .A1(program_cntr_out[6]), .A2(n431), .B1(N421), .B2(n154), 
        .ZN(n329) );
  INV_X1 U271 ( .A(n328), .ZN(n573) );
  AOI22_X1 U272 ( .A1(program_cntr_out[7]), .A2(n431), .B1(N422), .B2(n154), 
        .ZN(n328) );
  INV_X1 U273 ( .A(n327), .ZN(n572) );
  AOI22_X1 U274 ( .A1(program_cntr_out[8]), .A2(n212), .B1(N423), .B2(n154), 
        .ZN(n327) );
  INV_X1 U275 ( .A(n326), .ZN(n571) );
  AOI22_X1 U276 ( .A1(program_cntr_out[9]), .A2(n212), .B1(N424), .B2(n154), 
        .ZN(n326) );
  INV_X1 U277 ( .A(n325), .ZN(n570) );
  AOI22_X1 U278 ( .A1(program_cntr_out[10]), .A2(n212), .B1(N425), .B2(n154), 
        .ZN(n325) );
  INV_X1 U279 ( .A(n324), .ZN(n569) );
  AOI22_X1 U280 ( .A1(program_cntr_out[11]), .A2(n212), .B1(N426), .B2(n154), 
        .ZN(n324) );
  INV_X1 U281 ( .A(n323), .ZN(n568) );
  AOI22_X1 U282 ( .A1(program_cntr_out[12]), .A2(n187), .B1(N427), .B2(n155), 
        .ZN(n323) );
  INV_X1 U283 ( .A(n322), .ZN(n567) );
  AOI22_X1 U284 ( .A1(program_cntr_out[13]), .A2(n187), .B1(N428), .B2(n155), 
        .ZN(n322) );
  INV_X1 U285 ( .A(n321), .ZN(n566) );
  AOI22_X1 U286 ( .A1(program_cntr_out[14]), .A2(n187), .B1(N429), .B2(n155), 
        .ZN(n321) );
  INV_X1 U287 ( .A(n320), .ZN(n565) );
  AOI22_X1 U288 ( .A1(program_cntr_out[15]), .A2(n187), .B1(N430), .B2(n155), 
        .ZN(n320) );
  INV_X1 U289 ( .A(n319), .ZN(n564) );
  AOI22_X1 U290 ( .A1(program_cntr_out[16]), .A2(n186), .B1(N431), .B2(n155), 
        .ZN(n319) );
  INV_X1 U291 ( .A(n318), .ZN(n563) );
  AOI22_X1 U292 ( .A1(program_cntr_out[17]), .A2(n186), .B1(N432), .B2(n155), 
        .ZN(n318) );
  INV_X1 U293 ( .A(n377), .ZN(n622) );
  AOI22_X1 U294 ( .A1(initial_mask_out[22]), .A2(n443), .B1(N372), .B2(n151), 
        .ZN(n377) );
  INV_X1 U295 ( .A(n376), .ZN(n621) );
  AOI22_X1 U296 ( .A1(initial_mask_out[23]), .A2(n443), .B1(N373), .B2(n151), 
        .ZN(n376) );
  INV_X1 U297 ( .A(n375), .ZN(n620) );
  AOI22_X1 U298 ( .A1(initial_mask_out[24]), .A2(n443), .B1(N375), .B2(n151), 
        .ZN(n375) );
  INV_X1 U299 ( .A(n374), .ZN(n619) );
  AOI22_X1 U300 ( .A1(initial_mask_out[25]), .A2(n442), .B1(N376), .B2(n151), 
        .ZN(n374) );
  INV_X1 U301 ( .A(n373), .ZN(n618) );
  AOI22_X1 U302 ( .A1(initial_mask_out[26]), .A2(n442), .B1(N377), .B2(n151), 
        .ZN(n373) );
  INV_X1 U303 ( .A(n372), .ZN(n617) );
  AOI22_X1 U304 ( .A1(initial_mask_out[27]), .A2(n442), .B1(N378), .B2(n151), 
        .ZN(n372) );
  INV_X1 U305 ( .A(n371), .ZN(n616) );
  AOI22_X1 U306 ( .A1(initial_mask_out[28]), .A2(n442), .B1(N379), .B2(n151), 
        .ZN(n371) );
  INV_X1 U307 ( .A(n370), .ZN(n615) );
  AOI22_X1 U308 ( .A1(initial_mask_out[29]), .A2(n441), .B1(N380), .B2(n151), 
        .ZN(n370) );
  INV_X1 U309 ( .A(n369), .ZN(n614) );
  AOI22_X1 U310 ( .A1(initial_mask_out[30]), .A2(n441), .B1(N381), .B2(n151), 
        .ZN(n369) );
  INV_X1 U311 ( .A(n350), .ZN(n595) );
  AOI22_X1 U312 ( .A1(current_mask_out[17]), .A2(n436), .B1(N400), .B2(n153), 
        .ZN(n350) );
  INV_X1 U313 ( .A(n349), .ZN(n594) );
  AOI22_X1 U314 ( .A1(current_mask_out[18]), .A2(n436), .B1(N401), .B2(n153), 
        .ZN(n349) );
  INV_X1 U315 ( .A(n348), .ZN(n593) );
  AOI22_X1 U316 ( .A1(current_mask_out[19]), .A2(n436), .B1(N402), .B2(n153), 
        .ZN(n348) );
  INV_X1 U317 ( .A(n347), .ZN(n592) );
  AOI22_X1 U318 ( .A1(current_mask_out[20]), .A2(n436), .B1(N403), .B2(n153), 
        .ZN(n347) );
  INV_X1 U319 ( .A(n346), .ZN(n591) );
  AOI22_X1 U320 ( .A1(current_mask_out[21]), .A2(n435), .B1(N404), .B2(n153), 
        .ZN(n346) );
  INV_X1 U321 ( .A(n345), .ZN(n590) );
  AOI22_X1 U322 ( .A1(current_mask_out[22]), .A2(n435), .B1(N405), .B2(n153), 
        .ZN(n345) );
  INV_X1 U323 ( .A(n344), .ZN(n589) );
  AOI22_X1 U324 ( .A1(current_mask_out[23]), .A2(n435), .B1(N406), .B2(n153), 
        .ZN(n344) );
  INV_X1 U325 ( .A(n343), .ZN(n588) );
  AOI22_X1 U326 ( .A1(current_mask_out[24]), .A2(n435), .B1(N407), .B2(n153), 
        .ZN(n343) );
  INV_X1 U327 ( .A(n342), .ZN(n587) );
  AOI22_X1 U328 ( .A1(current_mask_out[25]), .A2(n434), .B1(N408), .B2(n153), 
        .ZN(n342) );
  INV_X1 U329 ( .A(n341), .ZN(n586) );
  AOI22_X1 U330 ( .A1(current_mask_out[26]), .A2(n434), .B1(N409), .B2(n151), 
        .ZN(n341) );
  INV_X1 U331 ( .A(n340), .ZN(n585) );
  AOI22_X1 U332 ( .A1(current_mask_out[27]), .A2(n434), .B1(N410), .B2(n154), 
        .ZN(n340) );
  INV_X1 U333 ( .A(n339), .ZN(n584) );
  AOI22_X1 U334 ( .A1(current_mask_out[28]), .A2(n434), .B1(N411), .B2(n154), 
        .ZN(n339) );
  INV_X1 U335 ( .A(n338), .ZN(n583) );
  AOI22_X1 U336 ( .A1(current_mask_out[29]), .A2(n433), .B1(N412), .B2(n151), 
        .ZN(n338) );
  INV_X1 U337 ( .A(n337), .ZN(n582) );
  AOI22_X1 U338 ( .A1(current_mask_out[30]), .A2(n433), .B1(N413), .B2(n153), 
        .ZN(n337) );
  INV_X1 U339 ( .A(n336), .ZN(n581) );
  AOI22_X1 U340 ( .A1(current_mask_out[31]), .A2(n433), .B1(N414), .B2(n151), 
        .ZN(n336) );
  INV_X1 U341 ( .A(n317), .ZN(n562) );
  AOI22_X1 U342 ( .A1(program_cntr_out[18]), .A2(n186), .B1(N433), .B2(n155), 
        .ZN(n317) );
  INV_X1 U343 ( .A(n316), .ZN(n561) );
  AOI22_X1 U344 ( .A1(program_cntr_out[19]), .A2(n186), .B1(N434), .B2(n155), 
        .ZN(n316) );
  INV_X1 U345 ( .A(n315), .ZN(n560) );
  AOI22_X1 U346 ( .A1(program_cntr_out[20]), .A2(n185), .B1(N435), .B2(n155), 
        .ZN(n315) );
  INV_X1 U347 ( .A(n314), .ZN(n559) );
  AOI22_X1 U348 ( .A1(program_cntr_out[21]), .A2(n185), .B1(N436), .B2(n156), 
        .ZN(n314) );
  INV_X1 U349 ( .A(n313), .ZN(n558) );
  AOI22_X1 U350 ( .A1(program_cntr_out[22]), .A2(n185), .B1(N437), .B2(n156), 
        .ZN(n313) );
  INV_X1 U351 ( .A(n312), .ZN(n557) );
  AOI22_X1 U352 ( .A1(program_cntr_out[23]), .A2(n185), .B1(N438), .B2(n156), 
        .ZN(n312) );
  INV_X1 U353 ( .A(n311), .ZN(n556) );
  AOI22_X1 U354 ( .A1(program_cntr_out[24]), .A2(n184), .B1(N439), .B2(n156), 
        .ZN(n311) );
  INV_X1 U355 ( .A(n310), .ZN(n555) );
  AOI22_X1 U356 ( .A1(program_cntr_out[25]), .A2(n184), .B1(N440), .B2(n156), 
        .ZN(n310) );
  INV_X1 U357 ( .A(n309), .ZN(n554) );
  AOI22_X1 U358 ( .A1(program_cntr_out[26]), .A2(n184), .B1(N441), .B2(n156), 
        .ZN(n309) );
  INV_X1 U359 ( .A(n308), .ZN(n553) );
  AOI22_X1 U360 ( .A1(program_cntr_out[27]), .A2(n184), .B1(N442), .B2(n156), 
        .ZN(n308) );
  INV_X1 U361 ( .A(n307), .ZN(n552) );
  AOI22_X1 U362 ( .A1(program_cntr_out[28]), .A2(n176), .B1(N443), .B2(n156), 
        .ZN(n307) );
  INV_X1 U363 ( .A(n306), .ZN(n551) );
  AOI22_X1 U364 ( .A1(program_cntr_out[29]), .A2(n176), .B1(N444), .B2(n156), 
        .ZN(n306) );
  INV_X1 U365 ( .A(n305), .ZN(n550) );
  AOI22_X1 U366 ( .A1(program_cntr_out[30]), .A2(n176), .B1(N445), .B2(n151), 
        .ZN(n305) );
  INV_X1 U367 ( .A(n246), .ZN(n499) );
  AOI22_X1 U368 ( .A1(n157), .A2(warp_lane_cnt[1]), .B1(n446), .B2(
        warp_lane_id_out[1]), .ZN(n246) );
  INV_X1 U369 ( .A(n236), .ZN(n498) );
  AOI22_X1 U370 ( .A1(n157), .A2(warp_lane_cnt[0]), .B1(n446), .B2(
        warp_lane_id_out[0]), .ZN(n236) );
  INV_X1 U371 ( .A(n218), .ZN(n497) );
  AOI22_X1 U372 ( .A1(n157), .A2(warp_id_cnt[1]), .B1(n446), .B2(
        warp_id_out[1]), .ZN(n218) );
  INV_X1 U373 ( .A(n304), .ZN(n549) );
  AOI22_X1 U374 ( .A1(program_cntr_out[31]), .A2(n176), .B1(N446), .B2(n154), 
        .ZN(n304) );
  INV_X1 U375 ( .A(n211), .ZN(n493) );
  AOI22_X1 U376 ( .A1(n152), .A2(warp_id_cnt[4]), .B1(n447), .B2(
        warp_id_out[4]), .ZN(n211) );
  INV_X1 U377 ( .A(n217), .ZN(n496) );
  AOI22_X1 U378 ( .A1(n157), .A2(warp_id_cnt[0]), .B1(n447), .B2(
        warp_id_out[0]), .ZN(n217) );
  INV_X1 U379 ( .A(n216), .ZN(n495) );
  AOI22_X1 U380 ( .A1(n152), .A2(warp_id_cnt[2]), .B1(n446), .B2(
        warp_id_out[2]), .ZN(n216) );
  INV_X1 U381 ( .A(n215), .ZN(n494) );
  AOI22_X1 U412 ( .A1(n157), .A2(warp_id_cnt[3]), .B1(n447), .B2(
        warp_id_out[3]), .ZN(n215) );
  INV_X1 U413 ( .A(n303), .ZN(n548) );
  AOI22_X1 U415 ( .A1(gprs_size_out[0]), .A2(n175), .B1(N447), .B2(n153), .ZN(
        n303) );
  INV_X1 U416 ( .A(n302), .ZN(n547) );
  AOI22_X1 U417 ( .A1(gprs_size_out[1]), .A2(n175), .B1(N448), .B2(n154), .ZN(
        n302) );
  INV_X1 U418 ( .A(n301), .ZN(n546) );
  AOI22_X1 U419 ( .A1(gprs_size_out[2]), .A2(n175), .B1(N449), .B2(n151), .ZN(
        n301) );
  INV_X1 U420 ( .A(n300), .ZN(n545) );
  AOI22_X1 U421 ( .A1(gprs_size_out[3]), .A2(n175), .B1(N450), .B2(n151), .ZN(
        n300) );
  INV_X1 U422 ( .A(n299), .ZN(n544) );
  AOI22_X1 U423 ( .A1(gprs_size_out[4]), .A2(n174), .B1(N451), .B2(n153), .ZN(
        n299) );
  INV_X1 U424 ( .A(n298), .ZN(n543) );
  AOI22_X1 U425 ( .A1(gprs_size_out[5]), .A2(n174), .B1(N452), .B2(n154), .ZN(
        n298) );
  INV_X1 U426 ( .A(n297), .ZN(n542) );
  AOI22_X1 U427 ( .A1(gprs_size_out[6]), .A2(n174), .B1(N453), .B2(n151), .ZN(
        n297) );
  INV_X1 U428 ( .A(n296), .ZN(n541) );
  AOI22_X1 U429 ( .A1(gprs_size_out[7]), .A2(n174), .B1(N454), .B2(n155), .ZN(
        n296) );
  INV_X1 U430 ( .A(n295), .ZN(n540) );
  AOI22_X1 U431 ( .A1(gprs_size_out[8]), .A2(n173), .B1(N455), .B2(n157), .ZN(
        n295) );
  INV_X1 U432 ( .A(n294), .ZN(n539) );
  AOI22_X1 U433 ( .A1(shmem_base_addr_out[0]), .A2(n173), .B1(N321), .B2(n156), 
        .ZN(n294) );
  INV_X1 U434 ( .A(n293), .ZN(n538) );
  AOI22_X1 U435 ( .A1(shmem_base_addr_out[1]), .A2(n173), .B1(N322), .B2(n152), 
        .ZN(n293) );
  INV_X1 U436 ( .A(n292), .ZN(n537) );
  AOI22_X1 U437 ( .A1(shmem_base_addr_out[2]), .A2(n173), .B1(N323), .B2(n153), 
        .ZN(n292) );
  INV_X1 U438 ( .A(n291), .ZN(n536) );
  AOI22_X1 U439 ( .A1(shmem_base_addr_out[3]), .A2(n172), .B1(N324), .B2(n153), 
        .ZN(n291) );
  INV_X1 U440 ( .A(n290), .ZN(n535) );
  AOI22_X1 U441 ( .A1(shmem_base_addr_out[4]), .A2(n172), .B1(N325), .B2(n155), 
        .ZN(n290) );
  INV_X1 U442 ( .A(n289), .ZN(n534) );
  AOI22_X1 U443 ( .A1(shmem_base_addr_out[5]), .A2(n172), .B1(N326), .B2(n157), 
        .ZN(n289) );
  INV_X1 U444 ( .A(n288), .ZN(n533) );
  AOI22_X1 U445 ( .A1(shmem_base_addr_out[6]), .A2(n172), .B1(N327), .B2(n156), 
        .ZN(n288) );
  INV_X1 U446 ( .A(n287), .ZN(n532) );
  AOI22_X1 U447 ( .A1(shmem_base_addr_out[7]), .A2(n171), .B1(N328), .B2(n151), 
        .ZN(n287) );
  INV_X1 U448 ( .A(n286), .ZN(n531) );
  AOI22_X1 U449 ( .A1(shmem_base_addr_out[8]), .A2(n171), .B1(N329), .B2(n152), 
        .ZN(n286) );
  INV_X1 U450 ( .A(n285), .ZN(n530) );
  AOI22_X1 U451 ( .A1(shmem_base_addr_out[9]), .A2(n431), .B1(N330), .B2(n153), 
        .ZN(n285) );
  INV_X1 U452 ( .A(n284), .ZN(n529) );
  AOI22_X1 U453 ( .A1(shmem_base_addr_out[10]), .A2(n171), .B1(N331), .B2(n154), .ZN(n284) );
  INV_X1 U454 ( .A(n283), .ZN(n528) );
  AOI22_X1 U455 ( .A1(shmem_base_addr_out[11]), .A2(n171), .B1(N332), .B2(n151), .ZN(n283) );
  INV_X1 U456 ( .A(n282), .ZN(n527) );
  AOI22_X1 U457 ( .A1(shmem_base_addr_out[12]), .A2(n165), .B1(N333), .B2(n152), .ZN(n282) );
  INV_X1 U458 ( .A(n281), .ZN(n526) );
  AOI22_X1 U459 ( .A1(shmem_base_addr_out[13]), .A2(n165), .B1(N334), .B2(n155), .ZN(n281) );
  INV_X1 U460 ( .A(n280), .ZN(n525) );
  AOI22_X1 U461 ( .A1(cta_id_out[0]), .A2(n165), .B1(N335), .B2(n156), .ZN(
        n280) );
  INV_X1 U462 ( .A(n279), .ZN(n524) );
  AOI22_X1 U463 ( .A1(cta_id_out[1]), .A2(n165), .B1(N336), .B2(n157), .ZN(
        n279) );
  INV_X1 U464 ( .A(n278), .ZN(n523) );
  AOI22_X1 U465 ( .A1(cta_id_out[2]), .A2(n164), .B1(N337), .B2(n151), .ZN(
        n278) );
  INV_X1 U466 ( .A(n277), .ZN(n522) );
  AOI22_X1 U467 ( .A1(cta_id_out[3]), .A2(n164), .B1(N338), .B2(n153), .ZN(
        n277) );
  INV_X1 U468 ( .A(n276), .ZN(n521) );
  AOI22_X1 U469 ( .A1(gprs_base_addr_out[0]), .A2(n164), .B1(N339), .B2(n153), 
        .ZN(n276) );
  INV_X1 U470 ( .A(n275), .ZN(n520) );
  AOI22_X1 U471 ( .A1(gprs_base_addr_out[1]), .A2(n164), .B1(N340), .B2(n151), 
        .ZN(n275) );
  INV_X1 U472 ( .A(n274), .ZN(n519) );
  AOI22_X1 U473 ( .A1(gprs_base_addr_out[2]), .A2(n163), .B1(N341), .B2(n154), 
        .ZN(n274) );
  INV_X1 U474 ( .A(n273), .ZN(n518) );
  AOI22_X1 U475 ( .A1(gprs_base_addr_out[3]), .A2(n163), .B1(N342), .B2(n154), 
        .ZN(n273) );
  INV_X1 U476 ( .A(n272), .ZN(n517) );
  AOI22_X1 U477 ( .A1(gprs_base_addr_out[4]), .A2(n163), .B1(N343), .B2(n154), 
        .ZN(n272) );
  INV_X1 U478 ( .A(n271), .ZN(n516) );
  AOI22_X1 U479 ( .A1(gprs_base_addr_out[5]), .A2(n163), .B1(N344), .B2(n154), 
        .ZN(n271) );
  INV_X1 U480 ( .A(n270), .ZN(n515) );
  AOI22_X1 U481 ( .A1(gprs_base_addr_out[6]), .A2(n162), .B1(N345), .B2(n153), 
        .ZN(n270) );
  INV_X1 U482 ( .A(n269), .ZN(n514) );
  AOI22_X1 U483 ( .A1(gprs_base_addr_out[7]), .A2(n162), .B1(N346), .B2(n155), 
        .ZN(n269) );
  INV_X1 U484 ( .A(n268), .ZN(n513) );
  AOI22_X1 U485 ( .A1(gprs_base_addr_out[8]), .A2(n162), .B1(N347), .B2(n155), 
        .ZN(n268) );
  INV_X1 U486 ( .A(n267), .ZN(n512) );
  AOI22_X1 U487 ( .A1(initial_mask_out[0]), .A2(n162), .B1(N348), .B2(n153), 
        .ZN(n267) );
  INV_X1 U488 ( .A(n266), .ZN(n511) );
  AOI22_X1 U489 ( .A1(initial_mask_out[1]), .A2(n160), .B1(N349), .B2(n153), 
        .ZN(n266) );
  INV_X1 U490 ( .A(n265), .ZN(n510) );
  AOI22_X1 U491 ( .A1(initial_mask_out[2]), .A2(n160), .B1(N350), .B2(n157), 
        .ZN(n265) );
  INV_X1 U492 ( .A(n264), .ZN(n509) );
  AOI22_X1 U493 ( .A1(initial_mask_out[3]), .A2(n160), .B1(N351), .B2(n156), 
        .ZN(n264) );
  INV_X1 U494 ( .A(n263), .ZN(n508) );
  AOI22_X1 U495 ( .A1(initial_mask_out[4]), .A2(n160), .B1(N352), .B2(n157), 
        .ZN(n263) );
  INV_X1 U496 ( .A(n262), .ZN(n507) );
  AOI22_X1 U497 ( .A1(initial_mask_out[5]), .A2(n159), .B1(N353), .B2(n155), 
        .ZN(n262) );
  INV_X1 U498 ( .A(n261), .ZN(n506) );
  AOI22_X1 U499 ( .A1(initial_mask_out[6]), .A2(n159), .B1(N354), .B2(n154), 
        .ZN(n261) );
  INV_X1 U500 ( .A(n386), .ZN(n631) );
  AOI22_X1 U501 ( .A1(initial_mask_out[13]), .A2(n445), .B1(N362), .B2(n156), 
        .ZN(n386) );
  INV_X1 U502 ( .A(n385), .ZN(n630) );
  AOI22_X1 U503 ( .A1(initial_mask_out[14]), .A2(n445), .B1(N364), .B2(n155), 
        .ZN(n385) );
  INV_X1 U504 ( .A(n384), .ZN(n629) );
  AOI22_X1 U505 ( .A1(initial_mask_out[15]), .A2(n445), .B1(N365), .B2(n153), 
        .ZN(n384) );
  INV_X1 U506 ( .A(n383), .ZN(n628) );
  AOI22_X1 U507 ( .A1(initial_mask_out[16]), .A2(n445), .B1(N366), .B2(n157), 
        .ZN(n383) );
  INV_X1 U508 ( .A(n382), .ZN(n627) );
  AOI22_X1 U509 ( .A1(initial_mask_out[17]), .A2(n444), .B1(N367), .B2(n152), 
        .ZN(n382) );
  INV_X1 U510 ( .A(n381), .ZN(n626) );
  AOI22_X1 U511 ( .A1(initial_mask_out[18]), .A2(n444), .B1(N368), .B2(n155), 
        .ZN(n381) );
  INV_X1 U512 ( .A(n380), .ZN(n625) );
  AOI22_X1 U513 ( .A1(initial_mask_out[19]), .A2(n444), .B1(N369), .B2(n156), 
        .ZN(n380) );
  INV_X1 U514 ( .A(n379), .ZN(n624) );
  AOI22_X1 U515 ( .A1(initial_mask_out[20]), .A2(n444), .B1(N370), .B2(n157), 
        .ZN(n379) );
  INV_X1 U516 ( .A(n378), .ZN(n623) );
  AOI22_X1 U517 ( .A1(initial_mask_out[21]), .A2(n443), .B1(N371), .B2(n157), 
        .ZN(n378) );
  INV_X1 U518 ( .A(n368), .ZN(n613) );
  AOI22_X1 U519 ( .A1(initial_mask_out[31]), .A2(n441), .B1(N382), .B2(n152), 
        .ZN(n368) );
  INV_X1 U520 ( .A(n367), .ZN(n612) );
  AOI22_X1 U521 ( .A1(current_mask_out[0]), .A2(n441), .B1(N383), .B2(n152), 
        .ZN(n367) );
  INV_X1 U522 ( .A(n366), .ZN(n611) );
  AOI22_X1 U523 ( .A1(current_mask_out[1]), .A2(n440), .B1(N384), .B2(n152), 
        .ZN(n366) );
  INV_X1 U524 ( .A(n365), .ZN(n610) );
  AOI22_X1 U525 ( .A1(current_mask_out[2]), .A2(n440), .B1(N385), .B2(n152), 
        .ZN(n365) );
  INV_X1 U526 ( .A(n364), .ZN(n609) );
  AOI22_X1 U527 ( .A1(current_mask_out[3]), .A2(n440), .B1(N386), .B2(n152), 
        .ZN(n364) );
  INV_X1 U528 ( .A(n363), .ZN(n608) );
  AOI22_X1 U529 ( .A1(current_mask_out[4]), .A2(n440), .B1(N387), .B2(n152), 
        .ZN(n363) );
  INV_X1 U530 ( .A(n362), .ZN(n607) );
  AOI22_X1 U531 ( .A1(current_mask_out[5]), .A2(n439), .B1(N388), .B2(n152), 
        .ZN(n362) );
  INV_X1 U532 ( .A(n361), .ZN(n606) );
  AOI22_X1 U533 ( .A1(current_mask_out[6]), .A2(n439), .B1(N389), .B2(n152), 
        .ZN(n361) );
  INV_X1 U534 ( .A(n360), .ZN(n605) );
  AOI22_X1 U535 ( .A1(current_mask_out[7]), .A2(n439), .B1(N390), .B2(n152), 
        .ZN(n360) );
  INV_X1 U536 ( .A(n359), .ZN(n604) );
  AOI22_X1 U537 ( .A1(current_mask_out[8]), .A2(n439), .B1(N391), .B2(n152), 
        .ZN(n359) );
  INV_X1 U538 ( .A(n358), .ZN(n603) );
  AOI22_X1 U539 ( .A1(current_mask_out[9]), .A2(n438), .B1(N392), .B2(n152), 
        .ZN(n358) );
  INV_X1 U540 ( .A(n357), .ZN(n602) );
  AOI22_X1 U541 ( .A1(current_mask_out[10]), .A2(n438), .B1(N393), .B2(n152), 
        .ZN(n357) );
  INV_X1 U542 ( .A(n356), .ZN(n601) );
  AOI22_X1 U543 ( .A1(current_mask_out[11]), .A2(n438), .B1(N394), .B2(n155), 
        .ZN(n356) );
  INV_X1 U544 ( .A(n355), .ZN(n600) );
  AOI22_X1 U545 ( .A1(current_mask_out[12]), .A2(n438), .B1(N395), .B2(n152), 
        .ZN(n355) );
  INV_X1 U546 ( .A(n354), .ZN(n599) );
  AOI22_X1 U547 ( .A1(current_mask_out[13]), .A2(n437), .B1(N396), .B2(n156), 
        .ZN(n354) );
  INV_X1 U548 ( .A(n353), .ZN(n598) );
  AOI22_X1 U549 ( .A1(current_mask_out[14]), .A2(n437), .B1(N397), .B2(n156), 
        .ZN(n353) );
  INV_X1 U550 ( .A(n352), .ZN(n597) );
  AOI22_X1 U551 ( .A1(current_mask_out[15]), .A2(n437), .B1(N398), .B2(n156), 
        .ZN(n352) );
  INV_X1 U552 ( .A(n351), .ZN(n596) );
  AOI22_X1 U553 ( .A1(current_mask_out[16]), .A2(n437), .B1(N399), .B2(n155), 
        .ZN(n351) );
  INV_X1 U554 ( .A(n260), .ZN(n505) );
  AOI22_X1 U555 ( .A1(initial_mask_out[7]), .A2(n159), .B1(N355), .B2(n157), 
        .ZN(n260) );
  INV_X1 U556 ( .A(n259), .ZN(n504) );
  AOI22_X1 U557 ( .A1(initial_mask_out[8]), .A2(n159), .B1(N356), .B2(n157), 
        .ZN(n259) );
  INV_X1 U558 ( .A(n258), .ZN(n503) );
  AOI22_X1 U559 ( .A1(initial_mask_out[9]), .A2(n158), .B1(N357), .B2(n157), 
        .ZN(n258) );
  INV_X1 U560 ( .A(n257), .ZN(n502) );
  AOI22_X1 U561 ( .A1(initial_mask_out[10]), .A2(n158), .B1(N358), .B2(n157), 
        .ZN(n257) );
  INV_X1 U562 ( .A(n256), .ZN(n501) );
  AOI22_X1 U563 ( .A1(initial_mask_out[11]), .A2(n158), .B1(N359), .B2(n157), 
        .ZN(n256) );
  INV_X1 U564 ( .A(n255), .ZN(n500) );
  AOI22_X1 U565 ( .A1(initial_mask_out[12]), .A2(n158), .B1(N360), .B2(n157), 
        .ZN(n255) );
  NOR3_X1 U566 ( .A1(n167), .A2(warp_scheduler_state_machine[1]), .A3(n161), 
        .ZN(n393) );
  OAI221_X1 U567 ( .B1(n188), .B2(n179), .C1(n632), .C2(n195), .A(n196), .ZN(
        n407) );
  OAI221_X1 U568 ( .B1(n188), .B2(n170), .C1(n632), .C2(n189), .A(n190), .ZN(
        n404) );
  OAI221_X1 U569 ( .B1(n188), .B2(n180), .C1(n632), .C2(n197), .A(n198), .ZN(
        n408) );
  OAI221_X1 U570 ( .B1(n188), .B2(n178), .C1(n632), .C2(n193), .A(n194), .ZN(
        n406) );
  OAI221_X1 U571 ( .B1(n188), .B2(n177), .C1(n632), .C2(n191), .A(n192), .ZN(
        n405) );
  OAI221_X1 U572 ( .B1(n639), .B2(n179), .C1(n202), .C2(n195), .A(n208), .ZN(
        n412) );
  OAI221_X1 U573 ( .B1(n639), .B2(n170), .C1(n202), .C2(n189), .A(n204), .ZN(
        n409) );
  OAI221_X1 U574 ( .B1(n639), .B2(n180), .C1(n202), .C2(n197), .A(n209), .ZN(
        n413) );
  OAI221_X1 U575 ( .B1(n639), .B2(n178), .C1(n202), .C2(n193), .A(n207), .ZN(
        n411) );
  OAI221_X1 U576 ( .B1(n639), .B2(n177), .C1(n202), .C2(n191), .A(n206), .ZN(
        n410) );
  NOR2_X1 U577 ( .A1(n168), .A2(n169), .ZN(n226) );
  OAI22_X1 U578 ( .A1(n161), .A2(n398), .B1(n490), .B2(n401), .ZN(n429) );
  AOI211_X1 U579 ( .C1(n393), .C2(warp_scheduler_next_state[2]), .A(n636), .B(
        n220), .ZN(n401) );
  OAI22_X1 U580 ( .A1(n167), .A2(n398), .B1(n490), .B2(n399), .ZN(n428) );
  AND3_X1 U581 ( .A1(n400), .A2(n639), .A3(n390), .ZN(n399) );
  AOI21_X1 U582 ( .B1(n393), .B2(warp_scheduler_next_state[0]), .A(n397), .ZN(
        n400) );
  OAI21_X1 U583 ( .B1(n390), .B2(pipeline_stall_in), .A(n640), .ZN(n389) );
  INV_X1 U584 ( .A(pipeline_stall_in), .ZN(n647) );
  OAI21_X1 U585 ( .B1(n227), .B2(n229), .A(n230), .ZN(n420) );
  AND3_X1 U586 ( .A1(n231), .A2(n131), .A3(n637), .ZN(n229) );
  OAI21_X1 U587 ( .B1(n131), .B2(n227), .A(n228), .ZN(n419) );
  OAI21_X1 U588 ( .B1(n387), .B2(n634), .A(n388), .ZN(n426) );
  INV_X1 U589 ( .A(n389), .ZN(n634) );
  NOR2_X1 U590 ( .A1(n245), .A2(n220), .ZN(n387) );
  OAI21_X1 U591 ( .B1(n240), .B2(n241), .A(n242), .ZN(n424) );
  AOI21_X1 U592 ( .B1(n243), .B2(n647), .A(n244), .ZN(n241) );
  NOR3_X1 U593 ( .A1(n225), .A2(n234), .A3(n245), .ZN(n240) );
  OAI21_X1 U594 ( .B1(n168), .B2(n237), .A(n247), .ZN(n425) );
  XNOR2_X1 U595 ( .A(n168), .B(warp_lane_cnt[0]), .ZN(n248) );
  OAI21_X1 U596 ( .B1(n169), .B2(n237), .A(n238), .ZN(n423) );
  INV_X1 U597 ( .A(n394), .ZN(n638) );
  AOI21_X1 U598 ( .B1(n392), .B2(done), .A(n395), .ZN(n394) );
  NOR3_X1 U599 ( .A1(n166), .A2(n167), .A3(n161), .ZN(n395) );
  NOR2_X1 U600 ( .A1(warp_state_rd_data_in[1]), .A2(warp_state_rd_data_in[0]), 
        .ZN(n254) );
  AND2_X1 U601 ( .A1(warp_state_rd_data_in[0]), .A2(warp_state_rd_data_in[1]), 
        .ZN(n219) );
  INV_X1 U602 ( .A(warp_state_rd_data_in[1]), .ZN(n649) );
  CLKBUF_X1 U603 ( .A(n134), .Z(n137) );
  CLKBUF_X1 U604 ( .A(n134), .Z(n138) );
  CLKBUF_X1 U605 ( .A(n134), .Z(n139) );
  CLKBUF_X1 U606 ( .A(n134), .Z(n140) );
  CLKBUF_X1 U607 ( .A(n134), .Z(n141) );
  CLKBUF_X1 U608 ( .A(n134), .Z(n142) );
  CLKBUF_X1 U609 ( .A(n135), .Z(n143) );
  CLKBUF_X1 U610 ( .A(n135), .Z(n144) );
  CLKBUF_X1 U611 ( .A(n135), .Z(n145) );
  CLKBUF_X1 U612 ( .A(n135), .Z(n146) );
  CLKBUF_X1 U613 ( .A(n135), .Z(n147) );
  CLKBUF_X1 U614 ( .A(n135), .Z(n148) );
  CLKBUF_X1 U615 ( .A(n136), .Z(n149) );
  CLKBUF_X1 U616 ( .A(n136), .Z(n150) );
  INV_X1 U617 ( .A(n448), .ZN(n151) );
  INV_X1 U618 ( .A(n448), .ZN(n153) );
  INV_X1 U619 ( .A(n449), .ZN(n155) );
  NOR2_X1 U620 ( .A1(num_warps_in[1]), .A2(num_warps_in[0]), .ZN(n464) );
  AOI21_X1 U621 ( .B1(num_warps_in[0]), .B2(num_warps_in[1]), .A(n464), .ZN(
        n463) );
  INV_X1 U622 ( .A(n463), .ZN(N63) );
  NAND2_X1 U623 ( .A1(n464), .A2(n467), .ZN(n465) );
  OAI21_X1 U624 ( .B1(n464), .B2(n467), .A(n465), .ZN(N64) );
  NOR2_X1 U625 ( .A1(num_warps_in[3]), .A2(n465), .ZN(n466) );
  XOR2_X1 U626 ( .A(num_warps_in[4]), .B(n466), .Z(N66) );
  XOR2_X1 U627 ( .A(\r149/carry[4] ), .B(warp_id_cnt[4]), .Z(N73) );
  NOR2_X1 U628 ( .A1(n178), .A2(N64), .ZN(n469) );
  NAND2_X1 U629 ( .A1(warp_id_cnt[3]), .A2(n133), .ZN(n481) );
  NOR2_X1 U630 ( .A1(n469), .A2(n487), .ZN(n472) );
  NAND2_X1 U631 ( .A1(warp_id_cnt[0]), .A2(num_warps_in[0]), .ZN(n468) );
  OAI21_X1 U632 ( .B1(n179), .B2(n468), .A(N63), .ZN(n470) );
  NAND2_X1 U633 ( .A1(N64), .A2(n178), .ZN(n478) );
  NOR2_X1 U634 ( .A1(n469), .A2(n486), .ZN(n475) );
  OAI211_X1 U635 ( .C1(warp_id_cnt[1]), .C2(n485), .A(n470), .B(n475), .ZN(
        n471) );
  NOR2_X1 U636 ( .A1(n133), .A2(warp_id_cnt[3]), .ZN(n477) );
  AOI21_X1 U637 ( .B1(n472), .B2(n471), .A(n477), .ZN(n473) );
  XNOR2_X1 U638 ( .A(warp_id_cnt[4]), .B(N66), .ZN(n480) );
  AOI22_X1 U639 ( .A1(n473), .A2(n480), .B1(warp_id_cnt[4]), .B2(n484), .ZN(
        N94) );
  NOR2_X1 U640 ( .A1(num_warps_in[0]), .A2(warp_id_cnt[0]), .ZN(n476) );
  AOI21_X1 U641 ( .B1(n179), .B2(n476), .A(N63), .ZN(n474) );
  OAI211_X1 U642 ( .C1(n476), .C2(n179), .A(n489), .B(n475), .ZN(n479) );
  NAND3_X1 U643 ( .A1(n479), .A2(n478), .A3(n488), .ZN(n482) );
  NAND3_X1 U644 ( .A1(n482), .A2(n481), .A3(n480), .ZN(n483) );
  OAI21_X1 U645 ( .B1(warp_id_cnt[4]), .B2(n484), .A(n483), .ZN(N67) );
endmodule
